clk_slow_inst : clk_slow PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
