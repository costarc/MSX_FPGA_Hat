library ieee ;
use ieee.std_logic_1164.all;

Entity C_74HC30 is
port (
	D: in std_logic_vector(7 downto 0);
	Y: out std_logic);
end C_74HC30;

Architecture behaviour of C_74HC30 is

	
begin

	Y  <= '0' when D = "11111111" else '1';
	
end behaviour;
