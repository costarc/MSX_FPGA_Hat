clock_25mhz_inst : clock_25mhz PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
