library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
	port(
		cs		: in std_logic;
		A		: in std_logic_vector(15 downto 0);
		D		: out std_logic_vector(7 downto 0)
	);
end rom;

architecture rtl of rom is
type ROM is array (0 to 32767) of std_logic_vector(7 downto 0);
constant galaga : rom := (
    x"41",
    x"42",
    x"17",
    x"40",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"07",
    x"47",
    x"41",
    x"4c",
    x"41",
    x"47",
    x"41",
    x"21",
    x"00",
    x"e0",
    x"11",
    x"01",
    x"e0",
    x"01",
    x"fe",
    x"0f",
    x"36",
    x"00",
    x"ed",
    x"b0",
    x"31",
    x"00",
    x"e7",
    x"cd",
    x"38",
    x"01",
    x"e6",
    x"cf",
    x"4f",
    x"e6",
    x"0c",
    x"87",
    x"87",
    x"b1",
    x"cd",
    x"3b",
    x"01",
    x"cd",
    x"ad",
    x"59",
    x"3e",
    x"c3",
    x"21",
    x"4c",
    x"40",
    x"32",
    x"9a",
    x"fd",
    x"22",
    x"9b",
    x"fd",
    x"fb",
    x"01",
    x"01",
    x"e2",
    x"cd",
    x"47",
    x"00",
    x"18",
    x"fe",
    x"31",
    x"00",
    x"e7",
    x"cd",
    x"3e",
    x"01",
    x"01",
    x"01",
    x"c2",
    x"cd",
    x"47",
    x"00",
    x"2a",
    x"09",
    x"e0",
    x"23",
    x"22",
    x"09",
    x"e0",
    x"cb",
    x"45",
    x"28",
    x"18",
    x"21",
    x"80",
    x"e7",
    x"f9",
    x"3e",
    x"20",
    x"5e",
    x"2c",
    x"56",
    x"2c",
    x"4e",
    x"2c",
    x"46",
    x"2c",
    x"c5",
    x"d5",
    x"3d",
    x"20",
    x"f3",
    x"21",
    x"00",
    x"e7",
    x"18",
    x"03",
    x"21",
    x"80",
    x"e7",
    x"11",
    x"00",
    x"1b",
    x"01",
    x"80",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"21",
    x"61",
    x"e0",
    x"7e",
    x"11",
    x"00",
    x"01",
    x"d5",
    x"cd",
    x"af",
    x"41",
    x"3a",
    x"60",
    x"e0",
    x"86",
    x"77",
    x"d1",
    x"cd",
    x"b3",
    x"41",
    x"23",
    x"7e",
    x"11",
    x"20",
    x"01",
    x"d5",
    x"cd",
    x"af",
    x"41",
    x"3a",
    x"60",
    x"e0",
    x"cb",
    x"2f",
    x"86",
    x"77",
    x"d1",
    x"cd",
    x"b3",
    x"41",
    x"cd",
    x"20",
    x"90",
    x"3e",
    x"0f",
    x"1e",
    x"8f",
    x"cd",
    x"93",
    x"00",
    x"3e",
    x"0e",
    x"cd",
    x"96",
    x"00",
    x"32",
    x"30",
    x"e0",
    x"3e",
    x"0f",
    x"1e",
    x"cf",
    x"cd",
    x"93",
    x"00",
    x"3e",
    x"0e",
    x"cd",
    x"96",
    x"00",
    x"21",
    x"30",
    x"e0",
    x"a6",
    x"77",
    x"3e",
    x"08",
    x"cd",
    x"41",
    x"01",
    x"32",
    x"31",
    x"e0",
    x"07",
    x"cb",
    x"11",
    x"07",
    x"07",
    x"07",
    x"cb",
    x"11",
    x"3a",
    x"30",
    x"e0",
    x"1f",
    x"1f",
    x"a1",
    x"f6",
    x"fc",
    x"2f",
    x"32",
    x"20",
    x"e0",
    x"3e",
    x"05",
    x"cd",
    x"41",
    x"01",
    x"32",
    x"32",
    x"e0",
    x"f6",
    x"5f",
    x"4f",
    x"0f",
    x"a1",
    x"0f",
    x"4f",
    x"3a",
    x"30",
    x"e0",
    x"a1",
    x"4f",
    x"87",
    x"a1",
    x"07",
    x"07",
    x"07",
    x"4f",
    x"3a",
    x"31",
    x"e0",
    x"a1",
    x"f6",
    x"fe",
    x"2f",
    x"21",
    x"22",
    x"e0",
    x"4e",
    x"77",
    x"47",
    x"79",
    x"2f",
    x"a0",
    x"32",
    x"21",
    x"e0",
    x"3e",
    x"06",
    x"cd",
    x"41",
    x"01",
    x"e6",
    x"02",
    x"3e",
    x"ff",
    x"28",
    x"02",
    x"3e",
    x"9c",
    x"08",
    x"3e",
    x"07",
    x"cd",
    x"41",
    x"01",
    x"4f",
    x"2f",
    x"47",
    x"3a",
    x"24",
    x"e0",
    x"a0",
    x"47",
    x"08",
    x"a0",
    x"32",
    x"23",
    x"e0",
    x"79",
    x"f6",
    x"00",
    x"32",
    x"24",
    x"e0",
    x"21",
    x"0c",
    x"e0",
    x"3a",
    x"23",
    x"e0",
    x"e6",
    x"10",
    x"28",
    x"04",
    x"7e",
    x"ee",
    x"01",
    x"77",
    x"7e",
    x"3d",
    x"ca",
    x"5a",
    x"41",
    x"11",
    x"00",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"3a",
    x"00",
    x"e0",
    x"3d",
    x"cc",
    x"29",
    x"86",
    x"c3",
    x"44",
    x"40",
    x"21",
    x"00",
    x"00",
    x"39",
    x"eb",
    x"f9",
    x"e1",
    x"d5",
    x"f9",
    x"c9",
    x"21",
    x"00",
    x"00",
    x"39",
    x"5d",
    x"54",
    x"7d",
    x"e6",
    x"e0",
    x"6f",
    x"f9",
    x"e1",
    x"d5",
    x"f9",
    x"c9",
    x"21",
    x"00",
    x"e5",
    x"11",
    x"97",
    x"41",
    x"06",
    x"0b",
    x"7d",
    x"c6",
    x"1e",
    x"77",
    x"2c",
    x"74",
    x"6f",
    x"1a",
    x"77",
    x"2c",
    x"13",
    x"1a",
    x"77",
    x"23",
    x"13",
    x"10",
    x"ef",
    x"c9",
    x"d7",
    x"41",
    x"35",
    x"46",
    x"04",
    x"4d",
    x"03",
    x"80",
    x"5a",
    x"87",
    x"4e",
    x"53",
    x"0b",
    x"57",
    x"e3",
    x"48",
    x"93",
    x"81",
    x"5e",
    x"5e",
    x"48",
    x"58",
    x"00",
    x"00",
    x"0e",
    x"00",
    x"18",
    x"02",
    x"0e",
    x"20",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"eb",
    x"79",
    x"cd",
    x"4d",
    x"00",
    x"7c",
    x"c6",
    x"08",
    x"67",
    x"79",
    x"cd",
    x"4d",
    x"00",
    x"7c",
    x"c6",
    x"08",
    x"67",
    x"79",
    x"cd",
    x"4d",
    x"00",
    x"eb",
    x"c9",
    x"cd",
    x"f4",
    x"88",
    x"cd",
    x"6e",
    x"41",
    x"3a",
    x"21",
    x"e0",
    x"a7",
    x"20",
    x"02",
    x"18",
    x"f5",
    x"cd",
    x"a1",
    x"8a",
    x"3e",
    x"01",
    x"32",
    x"00",
    x"e0",
    x"32",
    x"50",
    x"e2",
    x"32",
    x"58",
    x"e2",
    x"32",
    x"60",
    x"e2",
    x"cd",
    x"1e",
    x"5a",
    x"cd",
    x"e1",
    x"88",
    x"21",
    x"f8",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"cd",
    x"6e",
    x"41",
    x"cd",
    x"e5",
    x"85",
    x"3a",
    x"50",
    x"e2",
    x"a7",
    x"20",
    x"f4",
    x"21",
    x"f8",
    x"45",
    x"cd",
    x"8f",
    x"8a",
    x"21",
    x"05",
    x"46",
    x"cd",
    x"7e",
    x"8a",
    x"06",
    x"5a",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"c1",
    x"10",
    x"f9",
    x"cd",
    x"41",
    x"81",
    x"21",
    x"05",
    x"46",
    x"cd",
    x"8f",
    x"8a",
    x"cd",
    x"f7",
    x"5a",
    x"cd",
    x"79",
    x"5a",
    x"21",
    x"74",
    x"e0",
    x"36",
    x"ff",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"60",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"20",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"a0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"c0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"3a",
    x"74",
    x"e0",
    x"a7",
    x"20",
    x"d3",
    x"3a",
    x"0d",
    x"e0",
    x"fe",
    x"03",
    x"ca",
    x"f2",
    x"43",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"20",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"20",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"e0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"a0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"c0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"00",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"cd",
    x"e5",
    x"85",
    x"3a",
    x"28",
    x"e0",
    x"fe",
    x"03",
    x"ca",
    x"ec",
    x"42",
    x"fe",
    x"0b",
    x"ca",
    x"ec",
    x"42",
    x"fe",
    x"09",
    x"ca",
    x"ec",
    x"42",
    x"21",
    x"17",
    x"e0",
    x"7e",
    x"a7",
    x"28",
    x"32",
    x"34",
    x"47",
    x"3d",
    x"20",
    x"09",
    x"21",
    x"0d",
    x"e0",
    x"7e",
    x"32",
    x"19",
    x"e0",
    x"36",
    x"00",
    x"78",
    x"fe",
    x"78",
    x"da",
    x"e4",
    x"42",
    x"3e",
    x"78",
    x"32",
    x"17",
    x"e0",
    x"3a",
    x"d7",
    x"e4",
    x"a7",
    x"ca",
    x"0c",
    x"43",
    x"c3",
    x"6c",
    x"42",
    x"3a",
    x"28",
    x"e0",
    x"d6",
    x"0b",
    x"c2",
    x"6c",
    x"42",
    x"af",
    x"32",
    x"17",
    x"e0",
    x"c3",
    x"6c",
    x"42",
    x"3a",
    x"10",
    x"e0",
    x"21",
    x"d7",
    x"e4",
    x"b6",
    x"21",
    x"92",
    x"e0",
    x"b6",
    x"c2",
    x"6c",
    x"42",
    x"3a",
    x"28",
    x"e0",
    x"fe",
    x"05",
    x"ca",
    x"6c",
    x"42",
    x"c3",
    x"2c",
    x"42",
    x"af",
    x"32",
    x"17",
    x"e0",
    x"32",
    x"18",
    x"e0",
    x"3a",
    x"19",
    x"e0",
    x"32",
    x"0d",
    x"e0",
    x"3a",
    x"0e",
    x"e0",
    x"a7",
    x"ca",
    x"47",
    x"43",
    x"21",
    x"05",
    x"46",
    x"cd",
    x"7e",
    x"8a",
    x"06",
    x"5a",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"20",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"c1",
    x"10",
    x"ed",
    x"cd",
    x"41",
    x"81",
    x"21",
    x"05",
    x"46",
    x"cd",
    x"8f",
    x"8a",
    x"c3",
    x"6c",
    x"42",
    x"21",
    x"0f",
    x"46",
    x"cd",
    x"7e",
    x"8a",
    x"06",
    x"f0",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"20",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"c1",
    x"10",
    x"f3",
    x"cd",
    x"e5",
    x"89",
    x"cd",
    x"03",
    x"8a",
    x"21",
    x"b3",
    x"45",
    x"06",
    x"04",
    x"c5",
    x"cd",
    x"7e",
    x"8a",
    x"c1",
    x"10",
    x"f9",
    x"cd",
    x"36",
    x"8b",
    x"21",
    x"51",
    x"19",
    x"11",
    x"f6",
    x"e0",
    x"01",
    x"05",
    x"03",
    x"cd",
    x"4f",
    x"8a",
    x"21",
    x"b1",
    x"19",
    x"11",
    x"f9",
    x"e0",
    x"01",
    x"05",
    x"03",
    x"cd",
    x"4f",
    x"8a",
    x"2a",
    x"f0",
    x"e0",
    x"7c",
    x"b5",
    x"28",
    x"0a",
    x"2a",
    x"f2",
    x"e0",
    x"7c",
    x"b5",
    x"28",
    x"53",
    x"cd",
    x"59",
    x"8b",
    x"21",
    x"13",
    x"1a",
    x"11",
    x"fe",
    x"e0",
    x"01",
    x"01",
    x"02",
    x"cd",
    x"4f",
    x"8a",
    x"21",
    x"15",
    x"1a",
    x"3e",
    x"8d",
    x"cd",
    x"4d",
    x"00",
    x"21",
    x"17",
    x"1a",
    x"3e",
    x"6b",
    x"cd",
    x"4d",
    x"00",
    x"3e",
    x"01",
    x"32",
    x"c0",
    x"e2",
    x"32",
    x"c8",
    x"e2",
    x"32",
    x"d0",
    x"e2",
    x"01",
    x"00",
    x"06",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"c1",
    x"3a",
    x"21",
    x"e0",
    x"a7",
    x"20",
    x"05",
    x"0b",
    x"79",
    x"b0",
    x"20",
    x"f0",
    x"af",
    x"32",
    x"c0",
    x"e2",
    x"32",
    x"c8",
    x"e2",
    x"32",
    x"d0",
    x"e2",
    x"32",
    x"00",
    x"e0",
    x"cd",
    x"6e",
    x"41",
    x"cd",
    x"e5",
    x"89",
    x"c3",
    x"d7",
    x"41",
    x"21",
    x"ef",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"18",
    x"c4",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"e0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"a0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"c0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"00",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"cd",
    x"e5",
    x"85",
    x"3a",
    x"0d",
    x"e0",
    x"a7",
    x"c2",
    x"f2",
    x"43",
    x"21",
    x"59",
    x"44",
    x"af",
    x"f5",
    x"e5",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"a0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"c0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"cd",
    x"e5",
    x"85",
    x"e1",
    x"f1",
    x"be",
    x"3c",
    x"38",
    x"04",
    x"23",
    x"23",
    x"23",
    x"af",
    x"f5",
    x"e5",
    x"23",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"e9",
    x"96",
    x"a7",
    x"44",
    x"01",
    x"77",
    x"44",
    x"1e",
    x"a1",
    x"44",
    x"3c",
    x"aa",
    x"44",
    x"3c",
    x"b9",
    x"44",
    x"96",
    x"31",
    x"45",
    x"f0",
    x"fc",
    x"44",
    x"01",
    x"23",
    x"45",
    x"3c",
    x"a7",
    x"44",
    x"01",
    x"50",
    x"45",
    x"3a",
    x"a0",
    x"e0",
    x"fe",
    x"28",
    x"20",
    x"11",
    x"3e",
    x"01",
    x"32",
    x"88",
    x"e2",
    x"32",
    x"90",
    x"e2",
    x"32",
    x"98",
    x"e2",
    x"32",
    x"a3",
    x"e0",
    x"c3",
    x"29",
    x"44",
    x"3e",
    x"01",
    x"32",
    x"a0",
    x"e2",
    x"32",
    x"a8",
    x"e2",
    x"32",
    x"b8",
    x"e2",
    x"af",
    x"32",
    x"a3",
    x"e0",
    x"c3",
    x"29",
    x"44",
    x"21",
    x"6c",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"c3",
    x"29",
    x"44",
    x"21",
    x"13",
    x"19",
    x"11",
    x"a0",
    x"e0",
    x"01",
    x"01",
    x"01",
    x"cd",
    x"58",
    x"45",
    x"c3",
    x"29",
    x"44",
    x"3a",
    x"a3",
    x"e0",
    x"a7",
    x"21",
    x"8d",
    x"45",
    x"28",
    x"03",
    x"21",
    x"7d",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"21",
    x"a0",
    x"e0",
    x"7e",
    x"fe",
    x"28",
    x"20",
    x"02",
    x"36",
    x"64",
    x"cd",
    x"de",
    x"44",
    x"21",
    x"9b",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"c3",
    x"29",
    x"44",
    x"11",
    x"a0",
    x"e0",
    x"1a",
    x"fe",
    x"64",
    x"30",
    x"10",
    x"21",
    x"88",
    x"19",
    x"af",
    x"cd",
    x"4d",
    x"00",
    x"21",
    x"89",
    x"19",
    x"01",
    x"02",
    x"01",
    x"c3",
    x"58",
    x"45",
    x"21",
    x"95",
    x"45",
    x"c3",
    x"7e",
    x"8a",
    x"3a",
    x"b8",
    x"e2",
    x"a7",
    x"20",
    x"2f",
    x"3a",
    x"b0",
    x"e2",
    x"a7",
    x"20",
    x"08",
    x"3a",
    x"a3",
    x"e0",
    x"ee",
    x"01",
    x"32",
    x"b0",
    x"e2",
    x"21",
    x"a0",
    x"e0",
    x"7e",
    x"a7",
    x"28",
    x"10",
    x"35",
    x"11",
    x"00",
    x"01",
    x"cd",
    x"a4",
    x"85",
    x"cd",
    x"de",
    x"44",
    x"18",
    x"0e",
    x"af",
    x"08",
    x"18",
    x"10",
    x"af",
    x"32",
    x"b0",
    x"e2",
    x"21",
    x"a4",
    x"45",
    x"cd",
    x"8f",
    x"8a",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"10",
    x"08",
    x"3a",
    x"a3",
    x"e0",
    x"a7",
    x"ca",
    x"29",
    x"44",
    x"21",
    x"a7",
    x"45",
    x"08",
    x"20",
    x"06",
    x"cd",
    x"7e",
    x"8a",
    x"c3",
    x"29",
    x"44",
    x"cd",
    x"8f",
    x"8a",
    x"c3",
    x"29",
    x"44",
    x"cd",
    x"03",
    x"8a",
    x"e1",
    x"e1",
    x"c3",
    x"2c",
    x"42",
    x"c5",
    x"1a",
    x"11",
    x"30",
    x"e0",
    x"a7",
    x"28",
    x"07",
    x"47",
    x"af",
    x"c6",
    x"01",
    x"27",
    x"10",
    x"fb",
    x"12",
    x"c1",
    x"c3",
    x"4f",
    x"8a",
    x"04",
    x"19",
    x"0e",
    x"7e",
    x"85",
    x"7d",
    x"72",
    x"75",
    x"82",
    x"27",
    x"7f",
    x"76",
    x"20",
    x"78",
    x"79",
    x"84",
    x"83",
    x"46",
    x"19",
    x"0d",
    x"13",
    x"10",
    x"05",
    x"03",
    x"09",
    x"01",
    x"0c",
    x"22",
    x"02",
    x"0f",
    x"0e",
    x"15",
    x"13",
    x"4a",
    x"19",
    x"05",
    x"72",
    x"7f",
    x"7e",
    x"85",
    x"83",
    x"88",
    x"19",
    x"03",
    x"61",
    x"60",
    x"60",
    x"8b",
    x"19",
    x"06",
    x"60",
    x"60",
    x"00",
    x"80",
    x"84",
    x"83",
    x"8b",
    x"19",
    x"02",
    x"a9",
    x"18",
    x"09",
    x"10",
    x"05",
    x"12",
    x"06",
    x"05",
    x"03",
    x"14",
    x"27",
    x"1e",
    x"e8",
    x"18",
    x"09",
    x"1c",
    x"12",
    x"05",
    x"13",
    x"15",
    x"0c",
    x"14",
    x"13",
    x"1c",
    x"43",
    x"19",
    x"0b",
    x"83",
    x"78",
    x"7f",
    x"84",
    x"83",
    x"00",
    x"76",
    x"79",
    x"82",
    x"75",
    x"74",
    x"a3",
    x"19",
    x"0e",
    x"7e",
    x"85",
    x"7d",
    x"72",
    x"75",
    x"82",
    x"00",
    x"7f",
    x"76",
    x"00",
    x"78",
    x"79",
    x"84",
    x"83",
    x"03",
    x"1a",
    x"0e",
    x"78",
    x"79",
    x"84",
    x"8b",
    x"7d",
    x"79",
    x"83",
    x"83",
    x"00",
    x"82",
    x"71",
    x"84",
    x"79",
    x"7f",
    x"12",
    x"1a",
    x"06",
    x"61",
    x"60",
    x"60",
    x"8d",
    x"60",
    x"6b",
    x"68",
    x"19",
    x"0a",
    x"77",
    x"71",
    x"7d",
    x"75",
    x"00",
    x"83",
    x"84",
    x"71",
    x"82",
    x"84",
    x"a9",
    x"19",
    x"07",
    x"12",
    x"05",
    x"01",
    x"04",
    x"19",
    x"25",
    x"1e",
    x"a8",
    x"19",
    x"09",
    x"77",
    x"71",
    x"7d",
    x"75",
    x"00",
    x"7f",
    x"86",
    x"75",
    x"82",
    x"19",
    x"18",
    x"04",
    x"08",
    x"09",
    x"07",
    x"08",
    x"3a",
    x"18",
    x"05",
    x"13",
    x"03",
    x"0f",
    x"12",
    x"05",
    x"99",
    x"18",
    x"05",
    x"13",
    x"03",
    x"0f",
    x"12",
    x"05",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"d0",
    x"e8",
    x"06",
    x"0d",
    x"cd",
    x"e1",
    x"8a",
    x"21",
    x"51",
    x"e0",
    x"7e",
    x"3c",
    x"fe",
    x"09",
    x"38",
    x"0c",
    x"11",
    x"52",
    x"e0",
    x"1a",
    x"3c",
    x"fe",
    x"10",
    x"38",
    x"01",
    x"af",
    x"12",
    x"af",
    x"77",
    x"3d",
    x"fa",
    x"1e",
    x"47",
    x"87",
    x"87",
    x"87",
    x"21",
    x"78",
    x"48",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"e5",
    x"dd",
    x"e1",
    x"6e",
    x"26",
    x"ef",
    x"11",
    x"d0",
    x"e8",
    x"01",
    x"0c",
    x"00",
    x"ed",
    x"b0",
    x"0e",
    x"14",
    x"09",
    x"0e",
    x"0c",
    x"ed",
    x"b0",
    x"dd",
    x"7e",
    x"01",
    x"06",
    x"0c",
    x"12",
    x"1c",
    x"3c",
    x"3c",
    x"10",
    x"fa",
    x"06",
    x"0c",
    x"d6",
    x"17",
    x"12",
    x"1c",
    x"3c",
    x"3c",
    x"10",
    x"fa",
    x"3a",
    x"51",
    x"e0",
    x"3d",
    x"e6",
    x"06",
    x"21",
    x"89",
    x"e3",
    x"85",
    x"6f",
    x"4e",
    x"2c",
    x"46",
    x"ed",
    x"43",
    x"87",
    x"e3",
    x"79",
    x"ed",
    x"44",
    x"dd",
    x"86",
    x"07",
    x"4f",
    x"dd",
    x"7e",
    x"02",
    x"c6",
    x"5a",
    x"6f",
    x"26",
    x"e3",
    x"06",
    x"05",
    x"71",
    x"2c",
    x"10",
    x"fc",
    x"dd",
    x"6e",
    x"02",
    x"26",
    x"e3",
    x"7d",
    x"fe",
    x"19",
    x"08",
    x"3a",
    x"52",
    x"e0",
    x"4f",
    x"e6",
    x"07",
    x"cb",
    x"45",
    x"28",
    x"0f",
    x"11",
    x"c0",
    x"48",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"79",
    x"fe",
    x"08",
    x"38",
    x"0f",
    x"18",
    x"2b",
    x"11",
    x"c8",
    x"48",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"79",
    x"fe",
    x"08",
    x"38",
    x"1e",
    x"1a",
    x"eb",
    x"21",
    x"2d",
    x"00",
    x"19",
    x"07",
    x"4f",
    x"06",
    x"05",
    x"cb",
    x"01",
    x"30",
    x"02",
    x"35",
    x"35",
    x"1a",
    x"a7",
    x"28",
    x"03",
    x"cd",
    x"c8",
    x"47",
    x"13",
    x"23",
    x"10",
    x"ef",
    x"c3",
    x"41",
    x"48",
    x"1a",
    x"eb",
    x"21",
    x"2d",
    x"00",
    x"19",
    x"07",
    x"4f",
    x"06",
    x"05",
    x"cb",
    x"01",
    x"30",
    x"02",
    x"34",
    x"34",
    x"1a",
    x"a7",
    x"28",
    x"03",
    x"cd",
    x"c8",
    x"47",
    x"13",
    x"23",
    x"10",
    x"ef",
    x"c3",
    x"41",
    x"48",
    x"3a",
    x"53",
    x"e0",
    x"3c",
    x"32",
    x"53",
    x"e0",
    x"11",
    x"00",
    x"e3",
    x"21",
    x"49",
    x"18",
    x"06",
    x"04",
    x"c5",
    x"1a",
    x"13",
    x"d5",
    x"e5",
    x"3d",
    x"28",
    x"6b",
    x"3d",
    x"28",
    x"57",
    x"18",
    x"39",
    x"e1",
    x"d1",
    x"23",
    x"23",
    x"c1",
    x"10",
    x"ec",
    x"3a",
    x"52",
    x"e0",
    x"11",
    x"ff",
    x"ff",
    x"cb",
    x"5f",
    x"28",
    x"04",
    x"11",
    x"01",
    x"00",
    x"2f",
    x"e6",
    x"07",
    x"21",
    x"b8",
    x"48",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"4e",
    x"cb",
    x"41",
    x"28",
    x"07",
    x"2a",
    x"8f",
    x"e3",
    x"19",
    x"22",
    x"8f",
    x"e3",
    x"cb",
    x"49",
    x"28",
    x"07",
    x"2a",
    x"8d",
    x"e3",
    x"19",
    x"22",
    x"8d",
    x"e3",
    x"c3",
    x"32",
    x"46",
    x"e5",
    x"01",
    x"02",
    x"00",
    x"eb",
    x"6b",
    x"26",
    x"ef",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"11",
    x"20",
    x"00",
    x"19",
    x"eb",
    x"6b",
    x"26",
    x"ef",
    x"01",
    x"02",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"18",
    x"ab",
    x"eb",
    x"21",
    x"d0",
    x"48",
    x"3a",
    x"53",
    x"e0",
    x"e6",
    x"04",
    x"28",
    x"15",
    x"23",
    x"23",
    x"23",
    x"23",
    x"18",
    x"0f",
    x"eb",
    x"21",
    x"d8",
    x"48",
    x"3a",
    x"53",
    x"e0",
    x"e6",
    x"04",
    x"28",
    x"04",
    x"23",
    x"23",
    x"23",
    x"23",
    x"e5",
    x"d5",
    x"01",
    x"02",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"eb",
    x"e1",
    x"23",
    x"23",
    x"0e",
    x"02",
    x"cd",
    x"5c",
    x"00",
    x"c3",
    x"3a",
    x"47",
    x"7e",
    x"d9",
    x"d6",
    x"08",
    x"fe",
    x"60",
    x"38",
    x"02",
    x"d6",
    x"60",
    x"47",
    x"c5",
    x"06",
    x"00",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"4f",
    x"21",
    x"d0",
    x"e8",
    x"09",
    x"eb",
    x"21",
    x"18",
    x"00",
    x"19",
    x"0e",
    x"03",
    x"ed",
    x"b0",
    x"0e",
    x"09",
    x"eb",
    x"09",
    x"eb",
    x"09",
    x"0e",
    x"03",
    x"ed",
    x"b0",
    x"08",
    x"30",
    x"06",
    x"08",
    x"21",
    x"00",
    x"e9",
    x"18",
    x"04",
    x"08",
    x"21",
    x"00",
    x"ec",
    x"3a",
    x"52",
    x"e0",
    x"e6",
    x"02",
    x"20",
    x"04",
    x"01",
    x"80",
    x"01",
    x"09",
    x"ed",
    x"4b",
    x"87",
    x"e3",
    x"09",
    x"eb",
    x"c1",
    x"78",
    x"e6",
    x"07",
    x"4f",
    x"87",
    x"81",
    x"87",
    x"87",
    x"87",
    x"87",
    x"30",
    x"01",
    x"14",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"21",
    x"00",
    x"e8",
    x"78",
    x"e6",
    x"f8",
    x"87",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"06",
    x"10",
    x"1a",
    x"13",
    x"b6",
    x"77",
    x"23",
    x"10",
    x"f9",
    x"0e",
    x"20",
    x"eb",
    x"ed",
    x"b0",
    x"d9",
    x"c9",
    x"dd",
    x"e5",
    x"cd",
    x"6e",
    x"41",
    x"dd",
    x"e1",
    x"dd",
    x"5e",
    x"03",
    x"dd",
    x"56",
    x"04",
    x"21",
    x"00",
    x"e8",
    x"01",
    x"c0",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"dd",
    x"5e",
    x"05",
    x"dd",
    x"56",
    x"06",
    x"21",
    x"d0",
    x"e8",
    x"01",
    x"0c",
    x"00",
    x"e5",
    x"d5",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"eb",
    x"e1",
    x"0e",
    x"0c",
    x"09",
    x"cd",
    x"5c",
    x"00",
    x"c3",
    x"32",
    x"46",
    x"81",
    x"a0",
    x"05",
    x"00",
    x"05",
    x"81",
    x"18",
    x"1f",
    x"8d",
    x"b8",
    x"0a",
    x"c0",
    x"05",
    x"8d",
    x"18",
    x"1f",
    x"c1",
    x"d0",
    x"0f",
    x"80",
    x"06",
    x"c1",
    x"18",
    x"2f",
    x"cd",
    x"e8",
    x"14",
    x"40",
    x"07",
    x"cd",
    x"18",
    x"2f",
    x"01",
    x"a0",
    x"19",
    x"00",
    x"0d",
    x"01",
    x"19",
    x"3f",
    x"0d",
    x"b8",
    x"1e",
    x"c0",
    x"0d",
    x"0d",
    x"19",
    x"3f",
    x"41",
    x"d0",
    x"23",
    x"80",
    x"0e",
    x"41",
    x"19",
    x"4f",
    x"4d",
    x"e8",
    x"28",
    x"40",
    x"0f",
    x"4d",
    x"19",
    x"4f",
    x"00",
    x"01",
    x"03",
    x"01",
    x"03",
    x"00",
    x"03",
    x"01",
    x"70",
    x"60",
    x"58",
    x"60",
    x"74",
    x"48",
    x"70",
    x"60",
    x"1c",
    x"0c",
    x"34",
    x"0c",
    x"5c",
    x"24",
    x"1c",
    x"0c",
    x"90",
    x"92",
    x"91",
    x"93",
    x"94",
    x"96",
    x"95",
    x"97",
    x"98",
    x"9a",
    x"99",
    x"9b",
    x"9c",
    x"9e",
    x"9d",
    x"9f",
    x"cd",
    x"6e",
    x"41",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"20",
    x"f7",
    x"3a",
    x"0d",
    x"e0",
    x"e6",
    x"01",
    x"c2",
    x"70",
    x"4b",
    x"21",
    x"96",
    x"e0",
    x"7e",
    x"3d",
    x"c2",
    x"48",
    x"49",
    x"3a",
    x"10",
    x"e0",
    x"d6",
    x"05",
    x"fe",
    x"06",
    x"d2",
    x"48",
    x"49",
    x"34",
    x"21",
    x"2c",
    x"e3",
    x"06",
    x"28",
    x"7e",
    x"a7",
    x"20",
    x"0a",
    x"2d",
    x"10",
    x"f9",
    x"3c",
    x"32",
    x"96",
    x"e0",
    x"c3",
    x"48",
    x"49",
    x"3e",
    x"01",
    x"32",
    x"00",
    x"e2",
    x"45",
    x"36",
    x"00",
    x"0e",
    x"03",
    x"78",
    x"d6",
    x"05",
    x"38",
    x"03",
    x"0c",
    x"18",
    x"f9",
    x"cd",
    x"b0",
    x"4a",
    x"46",
    x"7d",
    x"e6",
    x"3c",
    x"87",
    x"87",
    x"6f",
    x"26",
    x"e4",
    x"36",
    x"05",
    x"2c",
    x"2c",
    x"ed",
    x"5b",
    x"98",
    x"e0",
    x"73",
    x"2c",
    x"72",
    x"7d",
    x"c6",
    x"08",
    x"6f",
    x"36",
    x"00",
    x"2c",
    x"70",
    x"3a",
    x"14",
    x"e0",
    x"a7",
    x"ca",
    x"01",
    x"4a",
    x"3a",
    x"8c",
    x"e0",
    x"a7",
    x"c2",
    x"01",
    x"4a",
    x"21",
    x"d7",
    x"e4",
    x"3a",
    x"8a",
    x"e0",
    x"3d",
    x"be",
    x"da",
    x"01",
    x"4a",
    x"21",
    x"8e",
    x"e0",
    x"34",
    x"3a",
    x"82",
    x"e0",
    x"3d",
    x"be",
    x"d2",
    x"01",
    x"4a",
    x"36",
    x"00",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"03",
    x"26",
    x"e3",
    x"6f",
    x"7e",
    x"a7",
    x"20",
    x"09",
    x"2d",
    x"f2",
    x"77",
    x"49",
    x"2e",
    x"03",
    x"c3",
    x"77",
    x"49",
    x"f5",
    x"e5",
    x"21",
    x"91",
    x"e0",
    x"7e",
    x"34",
    x"e1",
    x"4d",
    x"e6",
    x"01",
    x"47",
    x"3a",
    x"28",
    x"e0",
    x"a7",
    x"28",
    x"02",
    x"06",
    x"00",
    x"c5",
    x"78",
    x"87",
    x"45",
    x"21",
    x"13",
    x"4b",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"eb",
    x"78",
    x"a7",
    x"28",
    x"09",
    x"fe",
    x"03",
    x"28",
    x"03",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"01",
    x"4f",
    x"c6",
    x"04",
    x"08",
    x"d5",
    x"cd",
    x"b0",
    x"4a",
    x"7d",
    x"e6",
    x"3c",
    x"87",
    x"87",
    x"c6",
    x"0c",
    x"32",
    x"30",
    x"e0",
    x"d1",
    x"c1",
    x"f1",
    x"3d",
    x"28",
    x"02",
    x"36",
    x"04",
    x"05",
    x"ca",
    x"01",
    x"4a",
    x"79",
    x"c6",
    x"07",
    x"6f",
    x"26",
    x"e3",
    x"06",
    x"03",
    x"0e",
    x"02",
    x"7e",
    x"a7",
    x"28",
    x"10",
    x"c5",
    x"d5",
    x"e5",
    x"45",
    x"08",
    x"4f",
    x"08",
    x"cd",
    x"b0",
    x"4a",
    x"e1",
    x"d1",
    x"c1",
    x"0d",
    x"28",
    x"03",
    x"2c",
    x"10",
    x"e9",
    x"3a",
    x"30",
    x"e0",
    x"6f",
    x"26",
    x"e4",
    x"79",
    x"ed",
    x"44",
    x"c6",
    x"02",
    x"77",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"01",
    x"ca",
    x"46",
    x"4a",
    x"3a",
    x"15",
    x"e0",
    x"a7",
    x"ca",
    x"e0",
    x"48",
    x"21",
    x"8f",
    x"e0",
    x"34",
    x"3a",
    x"88",
    x"e0",
    x"be",
    x"d2",
    x"e0",
    x"48",
    x"36",
    x"00",
    x"cd",
    x"c2",
    x"8a",
    x"26",
    x"e3",
    x"e6",
    x"02",
    x"28",
    x"10",
    x"2e",
    x"0f",
    x"7e",
    x"a7",
    x"20",
    x"13",
    x"2c",
    x"7d",
    x"fe",
    x"19",
    x"38",
    x"f6",
    x"2e",
    x"05",
    x"18",
    x"f2",
    x"2e",
    x"18",
    x"7e",
    x"a7",
    x"20",
    x"03",
    x"2d",
    x"18",
    x"f9",
    x"45",
    x"cd",
    x"90",
    x"4a",
    x"c3",
    x"e0",
    x"48",
    x"3a",
    x"16",
    x"e0",
    x"a7",
    x"ca",
    x"e0",
    x"48",
    x"21",
    x"90",
    x"e0",
    x"34",
    x"3a",
    x"86",
    x"e0",
    x"be",
    x"d2",
    x"e0",
    x"48",
    x"36",
    x"00",
    x"cd",
    x"c2",
    x"8a",
    x"26",
    x"e3",
    x"cb",
    x"4f",
    x"28",
    x"04",
    x"2e",
    x"19",
    x"18",
    x"02",
    x"2e",
    x"23",
    x"e6",
    x"80",
    x"28",
    x"12",
    x"7e",
    x"a7",
    x"20",
    x"18",
    x"2c",
    x"7d",
    x"fe",
    x"2d",
    x"38",
    x"f6",
    x"2e",
    x"19",
    x"18",
    x"f2",
    x"7e",
    x"a7",
    x"20",
    x"0a",
    x"2d",
    x"7d",
    x"fe",
    x"19",
    x"30",
    x"f6",
    x"2e",
    x"2c",
    x"18",
    x"f2",
    x"45",
    x"cd",
    x"90",
    x"4a",
    x"c3",
    x"e0",
    x"48",
    x"0e",
    x"03",
    x"78",
    x"d6",
    x"05",
    x"38",
    x"03",
    x"0c",
    x"18",
    x"f9",
    x"79",
    x"fe",
    x"08",
    x"30",
    x"05",
    x"11",
    x"ec",
    x"8b",
    x"18",
    x"03",
    x"11",
    x"c8",
    x"8b",
    x"21",
    x"d7",
    x"e4",
    x"3a",
    x"8a",
    x"e0",
    x"3d",
    x"be",
    x"d8",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"21",
    x"00",
    x"e4",
    x"7e",
    x"a7",
    x"ca",
    x"c2",
    x"4a",
    x"7d",
    x"c6",
    x"10",
    x"6f",
    x"18",
    x"f5",
    x"af",
    x"cb",
    x"39",
    x"1f",
    x"cb",
    x"39",
    x"0c",
    x"0c",
    x"71",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"73",
    x"2c",
    x"72",
    x"2c",
    x"77",
    x"2c",
    x"2c",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"2c",
    x"70",
    x"2c",
    x"77",
    x"2c",
    x"3a",
    x"93",
    x"e0",
    x"77",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"36",
    x"00",
    x"11",
    x"12",
    x"e0",
    x"79",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"3d",
    x"12",
    x"7d",
    x"21",
    x"82",
    x"e7",
    x"e6",
    x"f0",
    x"0f",
    x"0f",
    x"85",
    x"6f",
    x"0d",
    x"79",
    x"0f",
    x"0f",
    x"0f",
    x"77",
    x"2c",
    x"11",
    x"58",
    x"e0",
    x"79",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"77",
    x"c9",
    x"2e",
    x"8c",
    x"18",
    x"8c",
    x"af",
    x"32",
    x"0d",
    x"e0",
    x"3e",
    x"03",
    x"32",
    x"a9",
    x"e0",
    x"c3",
    x"e0",
    x"48",
    x"3a",
    x"d7",
    x"e4",
    x"a7",
    x"c2",
    x"e0",
    x"48",
    x"23",
    x"7e",
    x"fe",
    x"fe",
    x"28",
    x"e7",
    x"fe",
    x"fc",
    x"28",
    x"0a",
    x"2a",
    x"d0",
    x"e4",
    x"11",
    x"06",
    x"00",
    x"19",
    x"22",
    x"d0",
    x"e4",
    x"21",
    x"00",
    x"e4",
    x"22",
    x"d2",
    x"e4",
    x"e6",
    x"01",
    x"47",
    x"3a",
    x"d5",
    x"e4",
    x"11",
    x"ae",
    x"4c",
    x"87",
    x"80",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"32",
    x"d6",
    x"e4",
    x"11",
    x"d8",
    x"e4",
    x"2a",
    x"d0",
    x"e4",
    x"7e",
    x"12",
    x"23",
    x"13",
    x"7e",
    x"12",
    x"23",
    x"22",
    x"d0",
    x"e4",
    x"d9",
    x"34",
    x"34",
    x"3e",
    x"08",
    x"32",
    x"a9",
    x"e0",
    x"21",
    x"d4",
    x"e4",
    x"7e",
    x"d9",
    x"47",
    x"2a",
    x"9e",
    x"e0",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"fe",
    x"ff",
    x"28",
    x"a0",
    x"4f",
    x"78",
    x"e6",
    x"01",
    x"11",
    x"d8",
    x"e4",
    x"83",
    x"5f",
    x"1a",
    x"47",
    x"11",
    x"dc",
    x"e4",
    x"1a",
    x"b8",
    x"30",
    x"05",
    x"3c",
    x"12",
    x"c3",
    x"e0",
    x"48",
    x"af",
    x"12",
    x"d9",
    x"34",
    x"d9",
    x"7e",
    x"47",
    x"23",
    x"fe",
    x"e8",
    x"30",
    x"15",
    x"fe",
    x"e0",
    x"38",
    x"2a",
    x"11",
    x"d6",
    x"e4",
    x"1a",
    x"3d",
    x"fa",
    x"9c",
    x"4b",
    x"12",
    x"78",
    x"e6",
    x"03",
    x"4f",
    x"06",
    x"ff",
    x"18",
    x"23",
    x"11",
    x"a8",
    x"e0",
    x"1a",
    x"3d",
    x"c2",
    x"70",
    x"4b",
    x"12",
    x"3c",
    x"32",
    x"a5",
    x"e0",
    x"21",
    x"c0",
    x"e4",
    x"22",
    x"d2",
    x"e4",
    x"0e",
    x"ff",
    x"06",
    x"04",
    x"18",
    x"0a",
    x"78",
    x"07",
    x"07",
    x"e6",
    x"03",
    x"4f",
    x"78",
    x"e6",
    x"3f",
    x"47",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"2a",
    x"d2",
    x"e4",
    x"79",
    x"3c",
    x"3c",
    x"77",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"ed",
    x"5b",
    x"d0",
    x"e4",
    x"3a",
    x"d4",
    x"e4",
    x"1f",
    x"30",
    x"03",
    x"13",
    x"13",
    x"13",
    x"1a",
    x"13",
    x"77",
    x"2c",
    x"1a",
    x"13",
    x"77",
    x"2c",
    x"1a",
    x"77",
    x"2c",
    x"2c",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"2c",
    x"70",
    x"2c",
    x"77",
    x"2c",
    x"36",
    x"01",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"2c",
    x"2c",
    x"22",
    x"d2",
    x"e4",
    x"7d",
    x"0f",
    x"0f",
    x"3d",
    x"21",
    x"80",
    x"e7",
    x"85",
    x"6f",
    x"11",
    x"58",
    x"e0",
    x"79",
    x"3c",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"77",
    x"c3",
    x"70",
    x"4b",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"b0",
    x"5f",
    x"80",
    x"b0",
    x"5f",
    x"00",
    x"08",
    x"00",
    x"b0",
    x"5f",
    x"80",
    x"b0",
    x"5f",
    x"00",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"08",
    x"b0",
    x"5f",
    x"00",
    x"b0",
    x"5f",
    x"00",
    x"08",
    x"08",
    x"b0",
    x"5f",
    x"80",
    x"b0",
    x"5f",
    x"80",
    x"08",
    x"08",
    x"c7",
    x"5f",
    x"80",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"08",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"9c",
    x"5f",
    x"00",
    x"b0",
    x"5f",
    x"00",
    x"08",
    x"00",
    x"9c",
    x"5f",
    x"80",
    x"b0",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"db",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"db",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"00",
    x"00",
    x"02",
    x"00",
    x"02",
    x"02",
    x"04",
    x"02",
    x"04",
    x"04",
    x"ff",
    x"fc",
    x"9d",
    x"49",
    x"9e",
    x"4a",
    x"e2",
    x"e1",
    x"a7",
    x"53",
    x"e2",
    x"e1",
    x"a8",
    x"54",
    x"ff",
    x"f1",
    x"00",
    x"48",
    x"e0",
    x"e1",
    x"01",
    x"4b",
    x"02",
    x"52",
    x"e0",
    x"e1",
    x"03",
    x"55",
    x"ff",
    x"f1",
    x"47",
    x"4c",
    x"e1",
    x"e1",
    x"46",
    x"4d",
    x"51",
    x"56",
    x"e1",
    x"e1",
    x"50",
    x"57",
    x"ff",
    x"f0",
    x"e2",
    x"e2",
    x"9c",
    x"9f",
    x"9b",
    x"a0",
    x"e2",
    x"e2",
    x"a6",
    x"a9",
    x"a5",
    x"aa",
    x"ff",
    x"f0",
    x"9a",
    x"a1",
    x"99",
    x"a2",
    x"a4",
    x"ab",
    x"e2",
    x"e2",
    x"e2",
    x"e2",
    x"a3",
    x"ac",
    x"e8",
    x"ff",
    x"fe",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"00",
    x"e4",
    x"dd",
    x"21",
    x"80",
    x"e7",
    x"06",
    x"0c",
    x"3a",
    x"a5",
    x"e0",
    x"a7",
    x"28",
    x"01",
    x"04",
    x"c5",
    x"e5",
    x"cd",
    x"28",
    x"4d",
    x"01",
    x"04",
    x"00",
    x"dd",
    x"09",
    x"e1",
    x"0e",
    x"10",
    x"09",
    x"c1",
    x"10",
    x"ef",
    x"c3",
    x"01",
    x"4d",
    x"e5",
    x"fd",
    x"e1",
    x"7e",
    x"a7",
    x"c8",
    x"3d",
    x"87",
    x"87",
    x"87",
    x"87",
    x"87",
    x"08",
    x"23",
    x"fd",
    x"7e",
    x"06",
    x"11",
    x"57",
    x"4d",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"47",
    x"7e",
    x"90",
    x"77",
    x"dc",
    x"5b",
    x"4d",
    x"23",
    x"23",
    x"23",
    x"7e",
    x"e6",
    x"7f",
    x"23",
    x"eb",
    x"21",
    x"12",
    x"4f",
    x"c3",
    x"f8",
    x"8a",
    x"04",
    x"07",
    x"0a",
    x"0e",
    x"23",
    x"5e",
    x"23",
    x"56",
    x"fd",
    x"35",
    x"0a",
    x"fa",
    x"66",
    x"4d",
    x"1b",
    x"1a",
    x"13",
    x"47",
    x"cb",
    x"7f",
    x"20",
    x"5b",
    x"23",
    x"4e",
    x"cb",
    x"09",
    x"cb",
    x"09",
    x"23",
    x"cb",
    x"77",
    x"20",
    x"1b",
    x"a9",
    x"cb",
    x"6f",
    x"7e",
    x"20",
    x"0a",
    x"3d",
    x"4f",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"0a",
    x"0d",
    x"18",
    x"07",
    x"3c",
    x"4f",
    x"e6",
    x"03",
    x"20",
    x"01",
    x"0c",
    x"79",
    x"e6",
    x"1f",
    x"77",
    x"2b",
    x"7e",
    x"e6",
    x"80",
    x"77",
    x"2b",
    x"72",
    x"2b",
    x"73",
    x"2b",
    x"78",
    x"e6",
    x"1f",
    x"87",
    x"87",
    x"86",
    x"77",
    x"f0",
    x"36",
    x"00",
    x"c9",
    x"e5",
    x"4d",
    x"ea",
    x"4d",
    x"ef",
    x"4d",
    x"fe",
    x"4d",
    x"06",
    x"4e",
    x"14",
    x"4e",
    x"32",
    x"4e",
    x"2b",
    x"4e",
    x"43",
    x"4e",
    x"4a",
    x"4e",
    x"63",
    x"4e",
    x"6d",
    x"4e",
    x"ad",
    x"4e",
    x"c1",
    x"4e",
    x"cf",
    x"4e",
    x"fb",
    x"4e",
    x"cb",
    x"77",
    x"20",
    x"09",
    x"e6",
    x"7f",
    x"e5",
    x"21",
    x"a8",
    x"4d",
    x"c3",
    x"f8",
    x"8a",
    x"e6",
    x"3f",
    x"fd",
    x"77",
    x"0a",
    x"18",
    x"8a",
    x"e1",
    x"72",
    x"2b",
    x"73",
    x"2b",
    x"c9",
    x"e1",
    x"18",
    x"81",
    x"fd",
    x"34",
    x"06",
    x"18",
    x"f8",
    x"fd",
    x"35",
    x"06",
    x"18",
    x"f3",
    x"1a",
    x"47",
    x"13",
    x"1a",
    x"13",
    x"fd",
    x"72",
    x"0f",
    x"fd",
    x"73",
    x"0e",
    x"57",
    x"58",
    x"18",
    x"e4",
    x"fd",
    x"56",
    x"0f",
    x"fd",
    x"5e",
    x"0e",
    x"18",
    x"dc",
    x"1a",
    x"13",
    x"47",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"b0",
    x"fd",
    x"77",
    x"04",
    x"18",
    x"c8",
    x"1a",
    x"47",
    x"13",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"20",
    x"05",
    x"fd",
    x"70",
    x"0d",
    x"18",
    x"bf",
    x"3e",
    x"1f",
    x"90",
    x"fd",
    x"77",
    x"0d",
    x"18",
    x"b7",
    x"1a",
    x"13",
    x"dd",
    x"77",
    x"00",
    x"18",
    x"b0",
    x"1a",
    x"13",
    x"fd",
    x"cb",
    x"04",
    x"7e",
    x"28",
    x"04",
    x"ed",
    x"44",
    x"c6",
    x"c0",
    x"dd",
    x"77",
    x"01",
    x"18",
    x"9f",
    x"1a",
    x"13",
    x"fd",
    x"77",
    x"06",
    x"18",
    x"98",
    x"1a",
    x"47",
    x"13",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"20",
    x"06",
    x"fd",
    x"70",
    x"05",
    x"c3",
    x"e2",
    x"4d",
    x"3e",
    x"1f",
    x"90",
    x"fd",
    x"77",
    x"05",
    x"c3",
    x"e2",
    x"4d",
    x"3a",
    x"dd",
    x"e4",
    x"a7",
    x"c2",
    x"e5",
    x"4d",
    x"c3",
    x"e2",
    x"4d",
    x"3a",
    x"93",
    x"e0",
    x"fd",
    x"77",
    x"0b",
    x"dd",
    x"e5",
    x"e1",
    x"7e",
    x"c6",
    x"30",
    x"77",
    x"3a",
    x"0d",
    x"e0",
    x"fe",
    x"02",
    x"20",
    x"1e",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"20",
    x"18",
    x"2c",
    x"7e",
    x"fd",
    x"cb",
    x"04",
    x"7e",
    x"28",
    x"04",
    x"ed",
    x"44",
    x"c6",
    x"c0",
    x"d6",
    x"70",
    x"f2",
    x"9a",
    x"4e",
    x"c6",
    x"50",
    x"c6",
    x"20",
    x"c3",
    x"34",
    x"4e",
    x"fd",
    x"7e",
    x"09",
    x"21",
    x"2d",
    x"e3",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"18",
    x"91",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"20",
    x"08",
    x"3a",
    x"0d",
    x"e0",
    x"fe",
    x"02",
    x"ca",
    x"e2",
    x"4d",
    x"11",
    x"ee",
    x"5f",
    x"c3",
    x"e2",
    x"4d",
    x"3a",
    x"85",
    x"e0",
    x"a7",
    x"ca",
    x"e2",
    x"4d",
    x"fd",
    x"36",
    x"06",
    x"02",
    x"c3",
    x"e2",
    x"4d",
    x"21",
    x"20",
    x"e1",
    x"7e",
    x"a7",
    x"c2",
    x"e2",
    x"4d",
    x"36",
    x"01",
    x"23",
    x"dd",
    x"7e",
    x"01",
    x"77",
    x"23",
    x"36",
    x"00",
    x"e1",
    x"e5",
    x"7d",
    x"e6",
    x"f0",
    x"32",
    x"25",
    x"e1",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"f6",
    x"09",
    x"fd",
    x"77",
    x"04",
    x"3e",
    x"01",
    x"32",
    x"b8",
    x"e1",
    x"c3",
    x"dc",
    x"4d",
    x"fd",
    x"7e",
    x"00",
    x"fe",
    x"02",
    x"ca",
    x"e2",
    x"4d",
    x"c3",
    x"fe",
    x"4d",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"c2",
    x"ef",
    x"4d",
    x"13",
    x"13",
    x"c3",
    x"e2",
    x"4d",
    x"34",
    x"4f",
    x"d9",
    x"4f",
    x"3f",
    x"50",
    x"c1",
    x"50",
    x"49",
    x"51",
    x"76",
    x"51",
    x"d5",
    x"4f",
    x"93",
    x"51",
    x"b6",
    x"51",
    x"94",
    x"52",
    x"83",
    x"51",
    x"ac",
    x"52",
    x"ce",
    x"51",
    x"fd",
    x"51",
    x"77",
    x"52",
    x"93",
    x"52",
    x"6e",
    x"51",
    x"eb",
    x"7e",
    x"47",
    x"23",
    x"7e",
    x"23",
    x"e6",
    x"03",
    x"28",
    x"5c",
    x"0f",
    x"0f",
    x"0f",
    x"80",
    x"11",
    x"80",
    x"9f",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"86",
    x"c6",
    x"08",
    x"47",
    x"fa",
    x"5a",
    x"4f",
    x"fe",
    x"10",
    x"38",
    x"10",
    x"e6",
    x"f0",
    x"18",
    x"02",
    x"f6",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"dd",
    x"86",
    x"00",
    x"dd",
    x"77",
    x"00",
    x"78",
    x"e6",
    x"0f",
    x"d6",
    x"08",
    x"77",
    x"23",
    x"7b",
    x"c6",
    x"08",
    x"e6",
    x"1f",
    x"47",
    x"7b",
    x"e6",
    x"e0",
    x"b0",
    x"5f",
    x"1a",
    x"86",
    x"c6",
    x"08",
    x"47",
    x"fa",
    x"88",
    x"4f",
    x"fe",
    x"10",
    x"38",
    x"10",
    x"e6",
    x"f0",
    x"18",
    x"02",
    x"f6",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"dd",
    x"86",
    x"01",
    x"dd",
    x"77",
    x"01",
    x"78",
    x"e6",
    x"0f",
    x"d6",
    x"08",
    x"77",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"7f",
    x"fe",
    x"02",
    x"28",
    x"0e",
    x"fd",
    x"7e",
    x"05",
    x"3c",
    x"3c",
    x"e6",
    x"1c",
    x"47",
    x"08",
    x"80",
    x"dd",
    x"77",
    x"02",
    x"c9",
    x"fd",
    x"7e",
    x"05",
    x"3c",
    x"3c",
    x"e6",
    x"1c",
    x"47",
    x"fd",
    x"be",
    x"0d",
    x"20",
    x"06",
    x"08",
    x"80",
    x"dd",
    x"77",
    x"02",
    x"c9",
    x"fd",
    x"7e",
    x"0d",
    x"e6",
    x"1c",
    x"b8",
    x"28",
    x"05",
    x"04",
    x"fd",
    x"70",
    x"0d",
    x"c9",
    x"fd",
    x"35",
    x"0d",
    x"c9",
    x"26",
    x"ff",
    x"18",
    x"02",
    x"26",
    x"00",
    x"fd",
    x"46",
    x"0d",
    x"78",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"05",
    x"78",
    x"3c",
    x"e6",
    x"1f",
    x"47",
    x"1a",
    x"4f",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"05",
    x"79",
    x"3c",
    x"e6",
    x"1f",
    x"4f",
    x"79",
    x"90",
    x"28",
    x"27",
    x"e6",
    x"1f",
    x"fe",
    x"10",
    x"30",
    x"0a",
    x"0d",
    x"79",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"0b",
    x"0d",
    x"18",
    x"08",
    x"0c",
    x"79",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"01",
    x"0c",
    x"79",
    x"e6",
    x"1f",
    x"12",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"24",
    x"ca",
    x"34",
    x"4f",
    x"c3",
    x"9a",
    x"4f",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"c9",
    x"06",
    x"04",
    x"11",
    x"ff",
    x"e2",
    x"13",
    x"1a",
    x"a7",
    x"20",
    x"02",
    x"10",
    x"f9",
    x"7b",
    x"32",
    x"a7",
    x"e0",
    x"87",
    x"87",
    x"87",
    x"87",
    x"c6",
    x"48",
    x"32",
    x"31",
    x"e3",
    x"c9",
    x"d5",
    x"fd",
    x"e5",
    x"e1",
    x"7e",
    x"3d",
    x"cc",
    x"25",
    x"50",
    x"fd",
    x"7e",
    x"09",
    x"fe",
    x"2d",
    x"30",
    x"52",
    x"c6",
    x"2d",
    x"6f",
    x"26",
    x"e3",
    x"5e",
    x"c6",
    x"2d",
    x"6f",
    x"56",
    x"dd",
    x"66",
    x"00",
    x"dd",
    x"6e",
    x"01",
    x"cd",
    x"d4",
    x"52",
    x"67",
    x"78",
    x"81",
    x"38",
    x"04",
    x"fe",
    x"08",
    x"38",
    x"2a",
    x"44",
    x"d1",
    x"1a",
    x"4f",
    x"90",
    x"28",
    x"18",
    x"e6",
    x"1f",
    x"fe",
    x"10",
    x"30",
    x"0a",
    x"0d",
    x"79",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"0b",
    x"0d",
    x"18",
    x"08",
    x"0c",
    x"79",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"01",
    x"0c",
    x"79",
    x"e6",
    x"1f",
    x"12",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"c3",
    x"34",
    x"4f",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"dd",
    x"72",
    x"00",
    x"dd",
    x"73",
    x"01",
    x"d1",
    x"c9",
    x"2c",
    x"36",
    x"00",
    x"11",
    x"b9",
    x"50",
    x"2c",
    x"73",
    x"2c",
    x"72",
    x"dd",
    x"56",
    x"00",
    x"dd",
    x"5e",
    x"01",
    x"cd",
    x"8a",
    x"59",
    x"fd",
    x"77",
    x"0d",
    x"d1",
    x"c9",
    x"88",
    x"02",
    x"84",
    x"06",
    x"cf",
    x"48",
    x"84",
    x"05",
    x"fd",
    x"7e",
    x"00",
    x"3d",
    x"28",
    x"46",
    x"fd",
    x"36",
    x"01",
    x"88",
    x"fd",
    x"34",
    x"04",
    x"13",
    x"13",
    x"af",
    x"12",
    x"26",
    x"e3",
    x"fd",
    x"7e",
    x"09",
    x"6f",
    x"fe",
    x"05",
    x"30",
    x"0b",
    x"dd",
    x"7e",
    x"03",
    x"fe",
    x"04",
    x"20",
    x"04",
    x"36",
    x"02",
    x"18",
    x"02",
    x"36",
    x"01",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"01",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"00",
    x"fd",
    x"7e",
    x"00",
    x"3d",
    x"3d",
    x"fe",
    x"03",
    x"28",
    x"3a",
    x"d0",
    x"21",
    x"14",
    x"e0",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"34",
    x"c9",
    x"fd",
    x"36",
    x"00",
    x"00",
    x"3e",
    x"05",
    x"32",
    x"28",
    x"e0",
    x"21",
    x"d7",
    x"e4",
    x"35",
    x"21",
    x"c0",
    x"e4",
    x"36",
    x"01",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"01",
    x"55",
    x"8c",
    x"71",
    x"2c",
    x"70",
    x"2c",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"80",
    x"77",
    x"7d",
    x"c6",
    x"06",
    x"6f",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"32",
    x"a5",
    x"e0",
    x"c9",
    x"fd",
    x"7e",
    x"09",
    x"21",
    x"15",
    x"e0",
    x"fe",
    x"19",
    x"38",
    x"01",
    x"23",
    x"34",
    x"c9",
    x"3a",
    x"51",
    x"e0",
    x"e6",
    x"01",
    x"c0",
    x"fd",
    x"7e",
    x"09",
    x"4f",
    x"26",
    x"e3",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"be",
    x"01",
    x"20",
    x"0b",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"be",
    x"00",
    x"20",
    x"01",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"c9",
    x"af",
    x"32",
    x"a5",
    x"e0",
    x"3c",
    x"32",
    x"a8",
    x"e0",
    x"21",
    x"d7",
    x"e4",
    x"35",
    x"fd",
    x"36",
    x"00",
    x"00",
    x"dd",
    x"36",
    x"00",
    x"e0",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"c0",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"f6",
    x"08",
    x"fd",
    x"77",
    x"04",
    x"18",
    x"07",
    x"fd",
    x"36",
    x"01",
    x"88",
    x"fd",
    x"34",
    x"04",
    x"fd",
    x"36",
    x"06",
    x"00",
    x"26",
    x"e3",
    x"fd",
    x"6e",
    x"09",
    x"36",
    x"00",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"01",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"00",
    x"c9",
    x"fd",
    x"7e",
    x"01",
    x"fe",
    x"09",
    x"d0",
    x"3e",
    x"01",
    x"32",
    x"08",
    x"e2",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"fd",
    x"77",
    x"04",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"f6",
    x"0d",
    x"fd",
    x"77",
    x"04",
    x"fd",
    x"36",
    x"06",
    x"00",
    x"26",
    x"e3",
    x"fd",
    x"7e",
    x"09",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"01",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"00",
    x"3e",
    x"3c",
    x"32",
    x"97",
    x"e0",
    x"fd",
    x"7e",
    x"09",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"21",
    x"97",
    x"e0",
    x"35",
    x"28",
    x"11",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"10",
    x"fd",
    x"7e",
    x"0c",
    x"20",
    x"03",
    x"3a",
    x"5c",
    x"e0",
    x"dd",
    x"77",
    x"03",
    x"c9",
    x"af",
    x"fd",
    x"77",
    x"01",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"fd",
    x"77",
    x"04",
    x"3a",
    x"5c",
    x"e0",
    x"dd",
    x"77",
    x"03",
    x"dd",
    x"36",
    x"02",
    x"80",
    x"eb",
    x"7d",
    x"e6",
    x"f0",
    x"6f",
    x"e5",
    x"11",
    x"a0",
    x"e4",
    x"01",
    x"10",
    x"00",
    x"ed",
    x"b0",
    x"e1",
    x"7d",
    x"0e",
    x"10",
    x"ed",
    x"b0",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"c6",
    x"80",
    x"6f",
    x"26",
    x"e7",
    x"e5",
    x"11",
    x"a8",
    x"e7",
    x"0e",
    x"04",
    x"ed",
    x"b0",
    x"e1",
    x"0e",
    x"04",
    x"ed",
    x"b0",
    x"3e",
    x"ff",
    x"32",
    x"a9",
    x"e4",
    x"32",
    x"b9",
    x"e4",
    x"2a",
    x"9a",
    x"e0",
    x"22",
    x"a2",
    x"e4",
    x"2a",
    x"9c",
    x"e0",
    x"22",
    x"b2",
    x"e4",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"34",
    x"3e",
    x"01",
    x"32",
    x"08",
    x"e2",
    x"c9",
    x"eb",
    x"2d",
    x"2d",
    x"56",
    x"2d",
    x"5e",
    x"2d",
    x"1a",
    x"87",
    x"87",
    x"77",
    x"2c",
    x"1a",
    x"13",
    x"73",
    x"2c",
    x"72",
    x"2c",
    x"2c",
    x"eb",
    x"fd",
    x"34",
    x"04",
    x"fd",
    x"36",
    x"06",
    x"00",
    x"c9",
    x"c9",
    x"3a",
    x"20",
    x"e1",
    x"a7",
    x"28",
    x"05",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"fd",
    x"77",
    x"04",
    x"c9",
    x"d5",
    x"eb",
    x"2d",
    x"2d",
    x"56",
    x"2d",
    x"5e",
    x"2d",
    x"36",
    x"7f",
    x"eb",
    x"dd",
    x"7e",
    x"00",
    x"96",
    x"f2",
    x"c0",
    x"52",
    x"ed",
    x"44",
    x"fe",
    x"04",
    x"d9",
    x"d1",
    x"d2",
    x"34",
    x"4f",
    x"d9",
    x"eb",
    x"36",
    x"00",
    x"2c",
    x"13",
    x"73",
    x"2c",
    x"72",
    x"d9",
    x"c3",
    x"34",
    x"4f",
    x"7c",
    x"c6",
    x"20",
    x"67",
    x"7a",
    x"c6",
    x"20",
    x"94",
    x"30",
    x"13",
    x"ed",
    x"44",
    x"4f",
    x"7b",
    x"95",
    x"30",
    x"07",
    x"ed",
    x"44",
    x"47",
    x"26",
    x"18",
    x"18",
    x"14",
    x"47",
    x"26",
    x"00",
    x"18",
    x"0f",
    x"4f",
    x"7b",
    x"95",
    x"30",
    x"07",
    x"ed",
    x"44",
    x"47",
    x"26",
    x"10",
    x"18",
    x"03",
    x"47",
    x"26",
    x"08",
    x"78",
    x"b9",
    x"38",
    x"06",
    x"41",
    x"4f",
    x"3e",
    x"04",
    x"84",
    x"67",
    x"79",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"6f",
    x"cb",
    x"3f",
    x"b8",
    x"30",
    x"0b",
    x"24",
    x"85",
    x"b8",
    x"30",
    x"06",
    x"24",
    x"87",
    x"b8",
    x"30",
    x"01",
    x"24",
    x"7c",
    x"21",
    x"2b",
    x"53",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"c9",
    x"00",
    x"01",
    x"02",
    x"04",
    x"08",
    x"06",
    x"05",
    x"04",
    x"10",
    x"0e",
    x"0d",
    x"0c",
    x"08",
    x"09",
    x"0a",
    x"0c",
    x"10",
    x"11",
    x"12",
    x"14",
    x"18",
    x"16",
    x"15",
    x"14",
    x"00",
    x"1e",
    x"1d",
    x"1c",
    x"18",
    x"19",
    x"1a",
    x"1c",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"57",
    x"53",
    x"3a",
    x"28",
    x"e0",
    x"c3",
    x"f8",
    x"8a",
    x"6f",
    x"53",
    x"ae",
    x"53",
    x"36",
    x"54",
    x"8e",
    x"55",
    x"34",
    x"56",
    x"80",
    x"56",
    x"6f",
    x"53",
    x"6f",
    x"53",
    x"04",
    x"54",
    x"58",
    x"55",
    x"03",
    x"55",
    x"e4",
    x"55",
    x"21",
    x"b4",
    x"e7",
    x"7e",
    x"fe",
    x"e0",
    x"28",
    x"d4",
    x"23",
    x"11",
    x"29",
    x"e0",
    x"3a",
    x"20",
    x"e0",
    x"a7",
    x"ca",
    x"4b",
    x"53",
    x"fe",
    x"03",
    x"ca",
    x"4b",
    x"53",
    x"0f",
    x"da",
    x"9c",
    x"53",
    x"7e",
    x"fe",
    x"b8",
    x"d2",
    x"4b",
    x"53",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"01",
    x"3c",
    x"86",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"7e",
    x"fe",
    x"08",
    x"da",
    x"4b",
    x"53",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"01",
    x"3d",
    x"3d",
    x"86",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"b5",
    x"e7",
    x"11",
    x"29",
    x"e0",
    x"3a",
    x"20",
    x"e0",
    x"a7",
    x"ca",
    x"4b",
    x"53",
    x"fe",
    x"03",
    x"ca",
    x"4b",
    x"53",
    x"0f",
    x"da",
    x"dc",
    x"53",
    x"7e",
    x"fe",
    x"aa",
    x"d2",
    x"4b",
    x"53",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"01",
    x"3c",
    x"86",
    x"77",
    x"2d",
    x"2d",
    x"2d",
    x"2d",
    x"c6",
    x"0d",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"7e",
    x"fe",
    x"08",
    x"da",
    x"4b",
    x"53",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"01",
    x"3d",
    x"3d",
    x"86",
    x"77",
    x"2d",
    x"2d",
    x"2d",
    x"2d",
    x"c6",
    x"0d",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"3e",
    x"08",
    x"32",
    x"28",
    x"e0",
    x"af",
    x"32",
    x"c0",
    x"e1",
    x"3a",
    x"63",
    x"e0",
    x"32",
    x"60",
    x"e0",
    x"21",
    x"b4",
    x"e7",
    x"34",
    x"7e",
    x"2c",
    x"2c",
    x"fe",
    x"a3",
    x"28",
    x"1b",
    x"11",
    x"29",
    x"e0",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"03",
    x"c2",
    x"4b",
    x"53",
    x"7e",
    x"a7",
    x"ca",
    x"4b",
    x"53",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"2c",
    x"36",
    x"0f",
    x"c3",
    x"4b",
    x"53",
    x"36",
    x"00",
    x"af",
    x"32",
    x"28",
    x"e0",
    x"32",
    x"18",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"c0",
    x"e1",
    x"7e",
    x"a7",
    x"20",
    x"01",
    x"34",
    x"af",
    x"32",
    x"b8",
    x"e1",
    x"3e",
    x"f0",
    x"32",
    x"60",
    x"e0",
    x"21",
    x"b4",
    x"e7",
    x"7e",
    x"fe",
    x"78",
    x"28",
    x"31",
    x"35",
    x"23",
    x"3a",
    x"21",
    x"e1",
    x"be",
    x"28",
    x"06",
    x"38",
    x"03",
    x"34",
    x"18",
    x"01",
    x"35",
    x"23",
    x"3a",
    x"25",
    x"e1",
    x"5f",
    x"16",
    x"e4",
    x"1a",
    x"a7",
    x"28",
    x"8d",
    x"11",
    x"29",
    x"e0",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"03",
    x"20",
    x"06",
    x"7e",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"21",
    x"22",
    x"e1",
    x"36",
    x"00",
    x"c3",
    x"4b",
    x"53",
    x"2c",
    x"2c",
    x"7e",
    x"a7",
    x"20",
    x"d8",
    x"21",
    x"20",
    x"e1",
    x"36",
    x"03",
    x"7d",
    x"c6",
    x"05",
    x"6f",
    x"7e",
    x"11",
    x"a6",
    x"e0",
    x"12",
    x"13",
    x"26",
    x"e4",
    x"3c",
    x"6f",
    x"36",
    x"00",
    x"2c",
    x"01",
    x"f8",
    x"5f",
    x"71",
    x"2c",
    x"70",
    x"2c",
    x"36",
    x"00",
    x"7d",
    x"c6",
    x"05",
    x"6f",
    x"7e",
    x"12",
    x"21",
    x"b4",
    x"e7",
    x"11",
    x"b0",
    x"e7",
    x"01",
    x"03",
    x"00",
    x"ed",
    x"b0",
    x"3e",
    x"08",
    x"12",
    x"13",
    x"3e",
    x"e0",
    x"12",
    x"21",
    x"28",
    x"e0",
    x"36",
    x"0a",
    x"af",
    x"32",
    x"c0",
    x"e1",
    x"32",
    x"29",
    x"e0",
    x"3c",
    x"21",
    x"c0",
    x"e4",
    x"77",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"01",
    x"55",
    x"8c",
    x"71",
    x"2c",
    x"70",
    x"2c",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"80",
    x"77",
    x"7d",
    x"c6",
    x"06",
    x"6f",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"21",
    x"f0",
    x"54",
    x"cd",
    x"7e",
    x"8a",
    x"c3",
    x"4b",
    x"53",
    x"85",
    x"19",
    x"10",
    x"76",
    x"79",
    x"77",
    x"78",
    x"84",
    x"75",
    x"82",
    x"00",
    x"73",
    x"71",
    x"80",
    x"84",
    x"85",
    x"82",
    x"75",
    x"74",
    x"21",
    x"29",
    x"e0",
    x"34",
    x"7e",
    x"fe",
    x"78",
    x"30",
    x"1b",
    x"fe",
    x"1e",
    x"20",
    x"0b",
    x"3e",
    x"01",
    x"32",
    x"38",
    x"e2",
    x"32",
    x"40",
    x"e2",
    x"32",
    x"48",
    x"e2",
    x"3a",
    x"a6",
    x"e0",
    x"6f",
    x"2c",
    x"26",
    x"e4",
    x"36",
    x"7f",
    x"c3",
    x"4b",
    x"53",
    x"3a",
    x"a6",
    x"e0",
    x"6f",
    x"2c",
    x"26",
    x"e4",
    x"36",
    x"00",
    x"21",
    x"f0",
    x"54",
    x"cd",
    x"8f",
    x"8a",
    x"3e",
    x"04",
    x"32",
    x"28",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"3e",
    x"09",
    x"32",
    x"28",
    x"e0",
    x"3e",
    x"01",
    x"32",
    x"18",
    x"e0",
    x"32",
    x"d8",
    x"e1",
    x"32",
    x"28",
    x"e2",
    x"32",
    x"30",
    x"e2",
    x"21",
    x"a5",
    x"e0",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"21",
    x"a6",
    x"e0",
    x"34",
    x"7e",
    x"fe",
    x"3c",
    x"38",
    x"09",
    x"3a",
    x"d7",
    x"e4",
    x"21",
    x"92",
    x"e0",
    x"b6",
    x"28",
    x"17",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"03",
    x"c2",
    x"7b",
    x"55",
    x"21",
    x"b2",
    x"e7",
    x"7e",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"2c",
    x"36",
    x"0f",
    x"c3",
    x"6f",
    x"53",
    x"3a",
    x"b4",
    x"e7",
    x"fe",
    x"e0",
    x"ca",
    x"df",
    x"55",
    x"3e",
    x"03",
    x"32",
    x"28",
    x"e0",
    x"21",
    x"b2",
    x"e7",
    x"7e",
    x"a7",
    x"28",
    x"0f",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"03",
    x"20",
    x"24",
    x"7e",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"18",
    x"1c",
    x"2d",
    x"7e",
    x"fe",
    x"67",
    x"28",
    x"08",
    x"38",
    x"03",
    x"35",
    x"18",
    x"11",
    x"34",
    x"18",
    x"0e",
    x"3a",
    x"b5",
    x"e7",
    x"fe",
    x"5a",
    x"20",
    x"07",
    x"2d",
    x"7e",
    x"fe",
    x"a3",
    x"28",
    x"14",
    x"34",
    x"21",
    x"b5",
    x"e7",
    x"7e",
    x"fe",
    x"5a",
    x"ca",
    x"4b",
    x"53",
    x"38",
    x"04",
    x"35",
    x"c3",
    x"4b",
    x"53",
    x"34",
    x"c3",
    x"4b",
    x"53",
    x"3e",
    x"01",
    x"32",
    x"28",
    x"e0",
    x"af",
    x"32",
    x"18",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"3e",
    x"0b",
    x"32",
    x"28",
    x"e0",
    x"21",
    x"b2",
    x"e7",
    x"7e",
    x"a7",
    x"28",
    x"11",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"03",
    x"c2",
    x"4b",
    x"53",
    x"7e",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"2d",
    x"7e",
    x"fe",
    x"60",
    x"28",
    x"0a",
    x"38",
    x"04",
    x"35",
    x"c3",
    x"4b",
    x"53",
    x"34",
    x"c3",
    x"4b",
    x"53",
    x"2d",
    x"7e",
    x"fe",
    x"a3",
    x"28",
    x"04",
    x"34",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"b0",
    x"e7",
    x"11",
    x"b4",
    x"e7",
    x"01",
    x"04",
    x"00",
    x"ed",
    x"b0",
    x"3e",
    x"e0",
    x"32",
    x"b0",
    x"e7",
    x"af",
    x"32",
    x"28",
    x"e0",
    x"32",
    x"17",
    x"e0",
    x"af",
    x"32",
    x"18",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"11",
    x"a7",
    x"e0",
    x"1a",
    x"6f",
    x"26",
    x"e3",
    x"7e",
    x"a7",
    x"c2",
    x"66",
    x"56",
    x"1b",
    x"1a",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"c6",
    x"80",
    x"6f",
    x"26",
    x"e7",
    x"11",
    x"b0",
    x"e7",
    x"7e",
    x"fe",
    x"68",
    x"f5",
    x"2c",
    x"c6",
    x"10",
    x"12",
    x"1c",
    x"7e",
    x"2c",
    x"12",
    x"f1",
    x"d2",
    x"4b",
    x"53",
    x"1c",
    x"7e",
    x"e6",
    x"1f",
    x"12",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"b0",
    x"e7",
    x"35",
    x"f2",
    x"4b",
    x"53",
    x"3e",
    x"01",
    x"32",
    x"17",
    x"e0",
    x"3e",
    x"05",
    x"32",
    x"28",
    x"e0",
    x"3a",
    x"63",
    x"e0",
    x"32",
    x"60",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"a7",
    x"e0",
    x"5e",
    x"4b",
    x"16",
    x"e3",
    x"eb",
    x"7e",
    x"a7",
    x"c2",
    x"6f",
    x"53",
    x"1b",
    x"1a",
    x"6f",
    x"26",
    x"e4",
    x"7e",
    x"fe",
    x"02",
    x"20",
    x"30",
    x"7d",
    x"c6",
    x"09",
    x"6f",
    x"7e",
    x"b9",
    x"20",
    x"28",
    x"af",
    x"32",
    x"a5",
    x"e0",
    x"1a",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"c6",
    x"80",
    x"6f",
    x"26",
    x"e7",
    x"11",
    x"b0",
    x"e7",
    x"7e",
    x"2c",
    x"d6",
    x"10",
    x"12",
    x"1c",
    x"7e",
    x"2c",
    x"12",
    x"1c",
    x"7e",
    x"e6",
    x"1f",
    x"12",
    x"c3",
    x"6f",
    x"53",
    x"7d",
    x"e6",
    x"f0",
    x"12",
    x"18",
    x"d8",
    x"21",
    x"00",
    x"e4",
    x"06",
    x"0c",
    x"7e",
    x"fe",
    x"02",
    x"28",
    x"08",
    x"7d",
    x"c6",
    x"10",
    x"6f",
    x"10",
    x"f5",
    x"18",
    x"0f",
    x"7d",
    x"c6",
    x"09",
    x"6f",
    x"7e",
    x"b9",
    x"ca",
    x"c1",
    x"56",
    x"7d",
    x"c6",
    x"07",
    x"6f",
    x"10",
    x"e4",
    x"21",
    x"b0",
    x"e7",
    x"7e",
    x"3c",
    x"c2",
    x"3e",
    x"55",
    x"2c",
    x"2c",
    x"7e",
    x"a7",
    x"c2",
    x"3e",
    x"55",
    x"3e",
    x"06",
    x"32",
    x"28",
    x"e0",
    x"3e",
    x"01",
    x"32",
    x"a5",
    x"e0",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"c3",
    x"6f",
    x"53",
    x"cd",
    x"6e",
    x"41",
    x"3a",
    x"b4",
    x"e7",
    x"d6",
    x"80",
    x"fe",
    x"28",
    x"d2",
    x"d3",
    x"57",
    x"3a",
    x"28",
    x"e0",
    x"fe",
    x"03",
    x"ca",
    x"d3",
    x"57",
    x"21",
    x"21",
    x"e0",
    x"7e",
    x"a7",
    x"20",
    x"10",
    x"23",
    x"7e",
    x"a7",
    x"ca",
    x"d3",
    x"57",
    x"21",
    x"25",
    x"e0",
    x"34",
    x"7e",
    x"fe",
    x"14",
    x"da",
    x"d3",
    x"57",
    x"af",
    x"32",
    x"25",
    x"e0",
    x"21",
    x"30",
    x"e1",
    x"11",
    x"06",
    x"00",
    x"06",
    x"02",
    x"cb",
    x"7e",
    x"28",
    x"06",
    x"19",
    x"10",
    x"f9",
    x"c3",
    x"d3",
    x"57",
    x"3e",
    x"01",
    x"32",
    x"90",
    x"e1",
    x"ed",
    x"5b",
    x"f0",
    x"e0",
    x"13",
    x"ed",
    x"53",
    x"f0",
    x"e0",
    x"3a",
    x"28",
    x"e0",
    x"3d",
    x"ca",
    x"aa",
    x"57",
    x"36",
    x"80",
    x"23",
    x"3a",
    x"b6",
    x"e7",
    x"4f",
    x"0f",
    x"11",
    x"9a",
    x"57",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"13",
    x"77",
    x"23",
    x"36",
    x"00",
    x"23",
    x"1a",
    x"77",
    x"23",
    x"36",
    x"00",
    x"21",
    x"b8",
    x"e7",
    x"05",
    x"20",
    x"04",
    x"7d",
    x"c6",
    x"04",
    x"6f",
    x"11",
    x"b4",
    x"e7",
    x"1a",
    x"1c",
    x"77",
    x"2c",
    x"1a",
    x"1c",
    x"77",
    x"2c",
    x"1a",
    x"c6",
    x"b0",
    x"77",
    x"2c",
    x"36",
    x"0f",
    x"c3",
    x"d3",
    x"57",
    x"b3",
    x"00",
    x"bf",
    x"41",
    x"00",
    x"4d",
    x"41",
    x"41",
    x"4d",
    x"00",
    x"41",
    x"bf",
    x"00",
    x"b3",
    x"bf",
    x"bf",
    x"36",
    x"81",
    x"23",
    x"36",
    x"b3",
    x"23",
    x"af",
    x"77",
    x"23",
    x"77",
    x"23",
    x"77",
    x"21",
    x"b8",
    x"e7",
    x"05",
    x"20",
    x"04",
    x"7d",
    x"c6",
    x"04",
    x"6f",
    x"11",
    x"b4",
    x"e7",
    x"1a",
    x"1c",
    x"77",
    x"2c",
    x"1a",
    x"1c",
    x"c6",
    x"06",
    x"77",
    x"2c",
    x"3e",
    x"d0",
    x"77",
    x"2c",
    x"36",
    x"0f",
    x"21",
    x"30",
    x"e1",
    x"11",
    x"b8",
    x"e7",
    x"06",
    x"02",
    x"e5",
    x"d5",
    x"cb",
    x"7e",
    x"ca",
    x"14",
    x"58",
    x"23",
    x"7e",
    x"23",
    x"cd",
    x"26",
    x"58",
    x"4f",
    x"1a",
    x"81",
    x"12",
    x"fe",
    x"f8",
    x"30",
    x"04",
    x"fe",
    x"b8",
    x"30",
    x"10",
    x"13",
    x"23",
    x"7e",
    x"23",
    x"cd",
    x"26",
    x"58",
    x"4f",
    x"1a",
    x"81",
    x"12",
    x"fe",
    x"ba",
    x"da",
    x"14",
    x"58",
    x"2a",
    x"f2",
    x"e0",
    x"23",
    x"22",
    x"f2",
    x"e0",
    x"3e",
    x"e0",
    x"d1",
    x"12",
    x"e1",
    x"36",
    x"00",
    x"18",
    x"02",
    x"d1",
    x"e1",
    x"7b",
    x"c6",
    x"04",
    x"5f",
    x"3e",
    x"06",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"10",
    x"b8",
    x"c3",
    x"08",
    x"57",
    x"86",
    x"fa",
    x"36",
    x"58",
    x"4f",
    x"e6",
    x"0f",
    x"77",
    x"79",
    x"e6",
    x"f0",
    x"1f",
    x"1f",
    x"1f",
    x"1f",
    x"c9",
    x"4f",
    x"f6",
    x"f0",
    x"77",
    x"79",
    x"2f",
    x"e6",
    x"f0",
    x"1f",
    x"1f",
    x"1f",
    x"1f",
    x"ed",
    x"44",
    x"c9",
    x"cd",
    x"6e",
    x"41",
    x"3a",
    x"0d",
    x"e0",
    x"3d",
    x"28",
    x"08",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"01",
    x"ca",
    x"fa",
    x"58",
    x"21",
    x"1a",
    x"e0",
    x"7e",
    x"a7",
    x"28",
    x"04",
    x"35",
    x"c3",
    x"fa",
    x"58",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"c2",
    x"fa",
    x"58",
    x"3a",
    x"80",
    x"e0",
    x"47",
    x"21",
    x"92",
    x"e0",
    x"7e",
    x"b8",
    x"d2",
    x"fa",
    x"58",
    x"21",
    x"a4",
    x"e0",
    x"7e",
    x"fe",
    x"30",
    x"38",
    x"02",
    x"3e",
    x"fc",
    x"c6",
    x"04",
    x"77",
    x"47",
    x"11",
    x"80",
    x"e7",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"3a",
    x"70",
    x"e0",
    x"e6",
    x"3c",
    x"0f",
    x"0f",
    x"c6",
    x"50",
    x"67",
    x"1a",
    x"bc",
    x"d2",
    x"fa",
    x"58",
    x"21",
    x"04",
    x"e4",
    x"78",
    x"87",
    x"87",
    x"85",
    x"6f",
    x"7e",
    x"e6",
    x"7f",
    x"c2",
    x"fa",
    x"58",
    x"2c",
    x"7e",
    x"97",
    x"fe",
    x"0b",
    x"30",
    x"4c",
    x"7d",
    x"c6",
    x"06",
    x"6f",
    x"7e",
    x"3d",
    x"fa",
    x"fa",
    x"58",
    x"77",
    x"21",
    x"92",
    x"e0",
    x"34",
    x"21",
    x"40",
    x"e1",
    x"7e",
    x"a7",
    x"28",
    x"06",
    x"2c",
    x"2c",
    x"2c",
    x"2c",
    x"18",
    x"f6",
    x"36",
    x"01",
    x"e5",
    x"01",
    x"80",
    x"06",
    x"09",
    x"1a",
    x"47",
    x"1c",
    x"77",
    x"2c",
    x"1a",
    x"4f",
    x"77",
    x"2c",
    x"e5",
    x"50",
    x"59",
    x"cd",
    x"8a",
    x"59",
    x"fe",
    x"12",
    x"20",
    x"02",
    x"3e",
    x"11",
    x"fe",
    x"00",
    x"20",
    x"02",
    x"3e",
    x"0e",
    x"4f",
    x"e1",
    x"36",
    x"c0",
    x"2c",
    x"36",
    x"0e",
    x"e1",
    x"2c",
    x"71",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"21",
    x"40",
    x"e1",
    x"dd",
    x"21",
    x"c0",
    x"e7",
    x"06",
    x"08",
    x"c5",
    x"7e",
    x"a7",
    x"28",
    x"05",
    x"e5",
    x"cd",
    x"19",
    x"59",
    x"e1",
    x"01",
    x"04",
    x"00",
    x"09",
    x"dd",
    x"09",
    x"c1",
    x"10",
    x"ed",
    x"c3",
    x"45",
    x"58",
    x"23",
    x"7e",
    x"4f",
    x"23",
    x"11",
    x"c0",
    x"9f",
    x"83",
    x"5f",
    x"1a",
    x"86",
    x"c6",
    x"08",
    x"47",
    x"fa",
    x"32",
    x"59",
    x"fe",
    x"10",
    x"38",
    x"15",
    x"e6",
    x"f0",
    x"18",
    x"02",
    x"f6",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"dd",
    x"86",
    x"00",
    x"fe",
    x"c0",
    x"d2",
    x"7d",
    x"59",
    x"dd",
    x"77",
    x"00",
    x"78",
    x"e6",
    x"0f",
    x"d6",
    x"08",
    x"77",
    x"23",
    x"7b",
    x"c6",
    x"08",
    x"e6",
    x"1f",
    x"47",
    x"7b",
    x"e6",
    x"e0",
    x"b0",
    x"5f",
    x"1a",
    x"86",
    x"c6",
    x"08",
    x"47",
    x"fa",
    x"65",
    x"59",
    x"fe",
    x"10",
    x"38",
    x"14",
    x"e6",
    x"f0",
    x"18",
    x"02",
    x"f6",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"dd",
    x"86",
    x"01",
    x"dd",
    x"77",
    x"01",
    x"fe",
    x"bc",
    x"30",
    x"07",
    x"78",
    x"e6",
    x"0f",
    x"d6",
    x"08",
    x"77",
    x"c9",
    x"2d",
    x"2d",
    x"2d",
    x"36",
    x"00",
    x"dd",
    x"36",
    x"00",
    x"e0",
    x"21",
    x"92",
    x"e0",
    x"35",
    x"c9",
    x"c5",
    x"21",
    x"b4",
    x"e7",
    x"7e",
    x"2c",
    x"6e",
    x"67",
    x"3a",
    x"28",
    x"e0",
    x"3d",
    x"20",
    x"04",
    x"7d",
    x"c6",
    x"07",
    x"6f",
    x"eb",
    x"cd",
    x"d4",
    x"52",
    x"c1",
    x"fe",
    x"0d",
    x"30",
    x"02",
    x"3e",
    x"0d",
    x"fe",
    x"13",
    x"d8",
    x"3e",
    x"12",
    x"c9",
    x"cd",
    x"a1",
    x"8a",
    x"cd",
    x"e5",
    x"89",
    x"cd",
    x"9c",
    x"95",
    x"cd",
    x"ae",
    x"98",
    x"cd",
    x"7d",
    x"41",
    x"cd",
    x"c4",
    x"59",
    x"21",
    x"02",
    x"e0",
    x"36",
    x"03",
    x"06",
    x"1e",
    x"cd",
    x"c2",
    x"8a",
    x"10",
    x"fb",
    x"21",
    x"01",
    x"ef",
    x"06",
    x"18",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"03",
    x"c6",
    x"20",
    x"cb",
    x"40",
    x"28",
    x"02",
    x"c6",
    x"04",
    x"77",
    x"2c",
    x"10",
    x"ef",
    x"21",
    x"01",
    x"ef",
    x"11",
    x"21",
    x"ef",
    x"06",
    x"df",
    x"c5",
    x"7e",
    x"a7",
    x"28",
    x"09",
    x"47",
    x"e6",
    x"fc",
    x"4f",
    x"04",
    x"78",
    x"e6",
    x"03",
    x"b1",
    x"12",
    x"1c",
    x"2c",
    x"c1",
    x"10",
    x"ec",
    x"06",
    x"18",
    x"cd",
    x"c2",
    x"8a",
    x"6f",
    x"e6",
    x"03",
    x"c6",
    x"03",
    x"4f",
    x"7d",
    x"e6",
    x"e0",
    x"80",
    x"6f",
    x"36",
    x"00",
    x"c6",
    x"20",
    x"6f",
    x"0d",
    x"20",
    x"f8",
    x"10",
    x"e8",
    x"21",
    x"01",
    x"ef",
    x"70",
    x"2c",
    x"70",
    x"c9",
    x"21",
    x"00",
    x"e1",
    x"06",
    x"01",
    x"cd",
    x"e1",
    x"8a",
    x"af",
    x"32",
    x"28",
    x"e0",
    x"32",
    x"a8",
    x"e0",
    x"af",
    x"32",
    x"45",
    x"e0",
    x"3e",
    x"03",
    x"32",
    x"47",
    x"e0",
    x"3e",
    x"07",
    x"32",
    x"48",
    x"e0",
    x"3e",
    x"ff",
    x"32",
    x"46",
    x"e0",
    x"21",
    x"40",
    x"e0",
    x"af",
    x"06",
    x"04",
    x"77",
    x"23",
    x"10",
    x"fc",
    x"3e",
    x"01",
    x"32",
    x"44",
    x"e0",
    x"01",
    x"00",
    x"00",
    x"ed",
    x"43",
    x"70",
    x"e0",
    x"ed",
    x"43",
    x"72",
    x"e0",
    x"af",
    x"32",
    x"75",
    x"e0",
    x"3e",
    x"03",
    x"32",
    x"0e",
    x"e0",
    x"cd",
    x"79",
    x"5a",
    x"cd",
    x"e8",
    x"5a",
    x"21",
    x"75",
    x"5a",
    x"11",
    x"58",
    x"e0",
    x"01",
    x"04",
    x"00",
    x"ed",
    x"b0",
    x"c9",
    x"06",
    x"0c",
    x"09",
    x"05",
    x"af",
    x"21",
    x"14",
    x"e0",
    x"77",
    x"23",
    x"77",
    x"23",
    x"77",
    x"21",
    x"30",
    x"e3",
    x"06",
    x"03",
    x"cd",
    x"e1",
    x"8a",
    x"11",
    x"2d",
    x"e3",
    x"21",
    x"dc",
    x"5a",
    x"01",
    x"04",
    x"00",
    x"ed",
    x"b0",
    x"21",
    x"32",
    x"e3",
    x"0e",
    x"04",
    x"3e",
    x"1d",
    x"06",
    x"0a",
    x"77",
    x"23",
    x"c6",
    x"0f",
    x"10",
    x"fa",
    x"0d",
    x"20",
    x"f3",
    x"3e",
    x"0f",
    x"06",
    x"04",
    x"21",
    x"5a",
    x"e3",
    x"77",
    x"23",
    x"10",
    x"fc",
    x"36",
    x"ff",
    x"21",
    x"51",
    x"e0",
    x"36",
    x"ff",
    x"23",
    x"36",
    x"00",
    x"21",
    x"10",
    x"e0",
    x"36",
    x"28",
    x"23",
    x"36",
    x"04",
    x"23",
    x"36",
    x"10",
    x"23",
    x"36",
    x"14",
    x"11",
    x"89",
    x"e3",
    x"21",
    x"e0",
    x"5a",
    x"0e",
    x"08",
    x"ed",
    x"b0",
    x"21",
    x"c0",
    x"e8",
    x"06",
    x"0c",
    x"c3",
    x"e1",
    x"8a",
    x"48",
    x"58",
    x"68",
    x"78",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"00",
    x"03",
    x"00",
    x"21",
    x"b0",
    x"e7",
    x"36",
    x"e0",
    x"23",
    x"36",
    x"75",
    x"23",
    x"36",
    x"00",
    x"23",
    x"36",
    x"0f",
    x"c9",
    x"af",
    x"32",
    x"d4",
    x"e4",
    x"32",
    x"dc",
    x"e4",
    x"32",
    x"d7",
    x"e4",
    x"32",
    x"91",
    x"e0",
    x"32",
    x"a0",
    x"e0",
    x"32",
    x"a1",
    x"e0",
    x"21",
    x"8c",
    x"e0",
    x"77",
    x"23",
    x"77",
    x"3c",
    x"32",
    x"0d",
    x"e0",
    x"21",
    x"8e",
    x"e0",
    x"77",
    x"2c",
    x"36",
    x"18",
    x"2c",
    x"36",
    x"20",
    x"21",
    x"75",
    x"e0",
    x"7e",
    x"4f",
    x"3c",
    x"fe",
    x"1b",
    x"38",
    x"02",
    x"3e",
    x"17",
    x"77",
    x"79",
    x"3c",
    x"3c",
    x"e6",
    x"03",
    x"ca",
    x"85",
    x"5c",
    x"79",
    x"3c",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"ed",
    x"44",
    x"81",
    x"87",
    x"4f",
    x"87",
    x"81",
    x"21",
    x"0d",
    x"5c",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"79",
    x"32",
    x"8b",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"4f",
    x"e6",
    x"0e",
    x"0f",
    x"eb",
    x"21",
    x"07",
    x"5c",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"22",
    x"d0",
    x"e4",
    x"eb",
    x"79",
    x"e6",
    x"01",
    x"32",
    x"dd",
    x"e4",
    x"78",
    x"32",
    x"d5",
    x"e4",
    x"cd",
    x"f7",
    x"5b",
    x"4f",
    x"87",
    x"81",
    x"32",
    x"87",
    x"e0",
    x"78",
    x"87",
    x"80",
    x"32",
    x"89",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"87",
    x"87",
    x"32",
    x"94",
    x"e0",
    x"78",
    x"87",
    x"80",
    x"32",
    x"83",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"4f",
    x"e6",
    x"08",
    x"32",
    x"85",
    x"e0",
    x"79",
    x"e6",
    x"07",
    x"32",
    x"23",
    x"e1",
    x"78",
    x"32",
    x"84",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"32",
    x"95",
    x"e0",
    x"78",
    x"32",
    x"96",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"32",
    x"aa",
    x"e0",
    x"78",
    x"32",
    x"60",
    x"e0",
    x"32",
    x"63",
    x"e0",
    x"3a",
    x"75",
    x"e0",
    x"3c",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"3d",
    x"fe",
    x"03",
    x"38",
    x"04",
    x"d6",
    x"03",
    x"18",
    x"f8",
    x"47",
    x"87",
    x"80",
    x"87",
    x"21",
    x"e5",
    x"5b",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"78",
    x"11",
    x"98",
    x"e0",
    x"01",
    x"06",
    x"00",
    x"ed",
    x"b0",
    x"cd",
    x"c6",
    x"95",
    x"21",
    x"b8",
    x"4c",
    x"22",
    x"9e",
    x"e0",
    x"c9",
    x"6d",
    x"8c",
    x"93",
    x"8c",
    x"96",
    x"8c",
    x"ab",
    x"8c",
    x"cf",
    x"8c",
    x"e2",
    x"8c",
    x"f2",
    x"8c",
    x"15",
    x"8d",
    x"2b",
    x"8d",
    x"7e",
    x"23",
    x"47",
    x"e6",
    x"f0",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"08",
    x"78",
    x"e6",
    x"0f",
    x"47",
    x"08",
    x"c9",
    x"36",
    x"4c",
    x"5e",
    x"4c",
    x"86",
    x"4c",
    x"40",
    x"00",
    x"00",
    x"46",
    x"00",
    x"04",
    x"80",
    x"11",
    x"00",
    x"47",
    x"20",
    x"04",
    x"01",
    x"21",
    x"11",
    x"37",
    x"21",
    x"b5",
    x"81",
    x"32",
    x"11",
    x"38",
    x"21",
    x"b5",
    x"41",
    x"42",
    x"21",
    x"38",
    x"21",
    x"b5",
    x"11",
    x"52",
    x"22",
    x"b9",
    x"21",
    x"d6",
    x"92",
    x"63",
    x"22",
    x"a9",
    x"31",
    x"d6",
    x"40",
    x"11",
    x"10",
    x"b7",
    x"01",
    x"d6",
    x"12",
    x"64",
    x"32",
    x"a7",
    x"31",
    x"e7",
    x"93",
    x"76",
    x"32",
    x"a8",
    x"41",
    x"e7",
    x"53",
    x"76",
    x"32",
    x"a8",
    x"41",
    x"e7",
    x"13",
    x"87",
    x"42",
    x"a9",
    x"41",
    x"b8",
    x"94",
    x"87",
    x"42",
    x"a9",
    x"61",
    x"b8",
    x"50",
    x"22",
    x"11",
    x"b7",
    x"21",
    x"b8",
    x"13",
    x"88",
    x"52",
    x"9a",
    x"61",
    x"d8",
    x"94",
    x"88",
    x"52",
    x"9a",
    x"61",
    x"d8",
    x"54",
    x"88",
    x"52",
    x"9c",
    x"61",
    x"d8",
    x"13",
    x"98",
    x"62",
    x"9c",
    x"71",
    x"e8",
    x"94",
    x"99",
    x"62",
    x"9c",
    x"71",
    x"e8",
    x"54",
    x"99",
    x"62",
    x"9c",
    x"71",
    x"e8",
    x"21",
    x"0d",
    x"e0",
    x"36",
    x"03",
    x"3e",
    x"1e",
    x"32",
    x"a2",
    x"e0",
    x"3a",
    x"71",
    x"e0",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"4f",
    x"e6",
    x"07",
    x"47",
    x"21",
    x"cf",
    x"5c",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"c5",
    x"cd",
    x"c6",
    x"95",
    x"c1",
    x"78",
    x"87",
    x"21",
    x"0b",
    x"5d",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"22",
    x"d0",
    x"e4",
    x"21",
    x"d7",
    x"5c",
    x"22",
    x"9e",
    x"e0",
    x"79",
    x"fe",
    x"06",
    x"3e",
    x"03",
    x"30",
    x"03",
    x"78",
    x"cb",
    x"3f",
    x"c6",
    x"0b",
    x"32",
    x"aa",
    x"e0",
    x"c9",
    x"05",
    x"06",
    x"03",
    x"00",
    x"07",
    x"01",
    x"02",
    x"04",
    x"ff",
    x"fc",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"ff",
    x"f1",
    x"c0",
    x"00",
    x"c0",
    x"00",
    x"c0",
    x"00",
    x"c0",
    x"00",
    x"ff",
    x"f1",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"ff",
    x"f0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"ff",
    x"f0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"ff",
    x"fe",
    x"1b",
    x"5d",
    x"43",
    x"5d",
    x"6b",
    x"5d",
    x"93",
    x"5d",
    x"bb",
    x"5d",
    x"e3",
    x"5d",
    x"0b",
    x"5e",
    x"33",
    x"5e",
    x"08",
    x"00",
    x"40",
    x"8d",
    x"00",
    x"40",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"52",
    x"8d",
    x"00",
    x"52",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"52",
    x"8d",
    x"80",
    x"52",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"40",
    x"8d",
    x"00",
    x"40",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"40",
    x"8d",
    x"80",
    x"40",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"6a",
    x"8d",
    x"00",
    x"6a",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"81",
    x"8d",
    x"00",
    x"81",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"81",
    x"8d",
    x"00",
    x"81",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"6a",
    x"8d",
    x"00",
    x"6a",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"6a",
    x"8d",
    x"80",
    x"6a",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"91",
    x"8d",
    x"00",
    x"a8",
    x"8d",
    x"00",
    x"08",
    x"00",
    x"bf",
    x"8d",
    x"00",
    x"bf",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"bf",
    x"8d",
    x"00",
    x"bf",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"91",
    x"8d",
    x"00",
    x"a8",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"91",
    x"8d",
    x"80",
    x"a8",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"e0",
    x"8d",
    x"00",
    x"db",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"fe",
    x"8d",
    x"00",
    x"fe",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"fe",
    x"8d",
    x"80",
    x"fe",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"e0",
    x"8d",
    x"00",
    x"db",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"db",
    x"8d",
    x"00",
    x"e0",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"2f",
    x"8e",
    x"00",
    x"2f",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"57",
    x"8e",
    x"00",
    x"57",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"57",
    x"8e",
    x"80",
    x"57",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"2f",
    x"8e",
    x"00",
    x"2f",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"2f",
    x"8e",
    x"80",
    x"2f",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"7a",
    x"8e",
    x"00",
    x"7a",
    x"8e",
    x"00",
    x"08",
    x"00",
    x"9f",
    x"8e",
    x"00",
    x"9f",
    x"8e",
    x"80",
    x"08",
    x"00",
    x"9f",
    x"8e",
    x"00",
    x"9f",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"7a",
    x"8e",
    x"00",
    x"7a",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"7a",
    x"8e",
    x"80",
    x"7a",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"bd",
    x"8e",
    x"00",
    x"bd",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"d9",
    x"8e",
    x"00",
    x"d9",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"d9",
    x"8e",
    x"80",
    x"d9",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"bd",
    x"8e",
    x"00",
    x"bd",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"bd",
    x"8e",
    x"80",
    x"bd",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"f5",
    x"8e",
    x"00",
    x"f5",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"09",
    x"8f",
    x"00",
    x"09",
    x"8f",
    x"00",
    x"08",
    x"08",
    x"09",
    x"8f",
    x"80",
    x"09",
    x"8f",
    x"80",
    x"08",
    x"08",
    x"f5",
    x"8e",
    x"00",
    x"f5",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"f5",
    x"8e",
    x"80",
    x"f5",
    x"8e",
    x"80",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"8c",
    x"e0",
    x"7e",
    x"3c",
    x"fe",
    x"3c",
    x"38",
    x"09",
    x"23",
    x"7e",
    x"3c",
    x"20",
    x"01",
    x"3d",
    x"77",
    x"af",
    x"2b",
    x"77",
    x"23",
    x"4e",
    x"79",
    x"06",
    x"00",
    x"fe",
    x"1e",
    x"38",
    x"06",
    x"04",
    x"fe",
    x"3c",
    x"38",
    x"01",
    x"04",
    x"11",
    x"87",
    x"e0",
    x"21",
    x"0f",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"11",
    x"89",
    x"e0",
    x"21",
    x"2d",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"79",
    x"06",
    x"00",
    x"fe",
    x"28",
    x"38",
    x"01",
    x"04",
    x"11",
    x"8b",
    x"e0",
    x"21",
    x"4b",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"3a",
    x"10",
    x"e0",
    x"06",
    x"00",
    x"fe",
    x"14",
    x"30",
    x"09",
    x"04",
    x"04",
    x"fe",
    x"0a",
    x"30",
    x"08",
    x"04",
    x"18",
    x"05",
    x"fe",
    x"1e",
    x"30",
    x"01",
    x"04",
    x"11",
    x"94",
    x"e0",
    x"21",
    x"73",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"3a",
    x"0d",
    x"e0",
    x"3d",
    x"3e",
    x"08",
    x"20",
    x"03",
    x"3a",
    x"95",
    x"e0",
    x"32",
    x"80",
    x"e0",
    x"05",
    x"f2",
    x"d7",
    x"5e",
    x"06",
    x"00",
    x"11",
    x"83",
    x"e0",
    x"21",
    x"93",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"3a",
    x"17",
    x"e0",
    x"a7",
    x"c2",
    x"5b",
    x"5e",
    x"21",
    x"10",
    x"e0",
    x"3a",
    x"84",
    x"e0",
    x"be",
    x"da",
    x"5b",
    x"5e",
    x"21",
    x"0d",
    x"e0",
    x"7e",
    x"3d",
    x"ca",
    x"5b",
    x"5e",
    x"3e",
    x"02",
    x"77",
    x"3e",
    x"07",
    x"32",
    x"8a",
    x"e0",
    x"c3",
    x"5b",
    x"5e",
    x"1a",
    x"80",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"1b",
    x"12",
    x"c9",
    x"60",
    x"50",
    x"40",
    x"50",
    x"40",
    x"30",
    x"50",
    x"30",
    x"30",
    x"40",
    x"30",
    x"20",
    x"40",
    x"20",
    x"20",
    x"30",
    x"30",
    x"20",
    x"30",
    x"20",
    x"10",
    x"20",
    x"20",
    x"10",
    x"20",
    x"10",
    x"10",
    x"10",
    x"10",
    x"10",
    x"90",
    x"70",
    x"50",
    x"80",
    x"60",
    x"40",
    x"70",
    x"50",
    x"40",
    x"60",
    x"40",
    x"30",
    x"50",
    x"30",
    x"30",
    x"40",
    x"30",
    x"30",
    x"40",
    x"20",
    x"20",
    x"30",
    x"30",
    x"20",
    x"30",
    x"20",
    x"20",
    x"20",
    x"20",
    x"20",
    x"02",
    x"02",
    x"02",
    x"03",
    x"02",
    x"03",
    x"02",
    x"03",
    x"03",
    x"03",
    x"03",
    x"03",
    x"03",
    x"04",
    x"02",
    x"03",
    x"03",
    x"04",
    x"04",
    x"04",
    x"04",
    x"05",
    x"04",
    x"05",
    x"04",
    x"05",
    x"02",
    x"03",
    x"04",
    x"06",
    x"05",
    x"06",
    x"05",
    x"06",
    x"05",
    x"07",
    x"05",
    x"07",
    x"05",
    x"07",
    x"01",
    x"01",
    x"02",
    x"02",
    x"01",
    x"02",
    x"02",
    x"02",
    x"01",
    x"02",
    x"02",
    x"03",
    x"02",
    x"02",
    x"02",
    x"03",
    x"02",
    x"02",
    x"03",
    x"03",
    x"02",
    x"02",
    x"03",
    x"04",
    x"02",
    x"03",
    x"03",
    x"04",
    x"03",
    x"03",
    x"03",
    x"04",
    x"07",
    x"05",
    x"03",
    x"06",
    x"04",
    x"02",
    x"05",
    x"03",
    x"02",
    x"89",
    x"08",
    x"86",
    x"08",
    x"87",
    x"70",
    x"88",
    x"02",
    x"03",
    x"03",
    x"c7",
    x"48",
    x"c9",
    x"04",
    x"8a",
    x"c8",
    x"04",
    x"82",
    x"ee",
    x"5f",
    x"89",
    x"08",
    x"86",
    x"08",
    x"87",
    x"80",
    x"88",
    x"02",
    x"03",
    x"03",
    x"58",
    x"58",
    x"80",
    x"58",
    x"c9",
    x"07",
    x"81",
    x"8a",
    x"c8",
    x"07",
    x"82",
    x"ee",
    x"5f",
    x"89",
    x"0f",
    x"86",
    x"50",
    x"87",
    x"f1",
    x"88",
    x"02",
    x"50",
    x"c2",
    x"06",
    x"0a",
    x"c4",
    x"50",
    x"8a",
    x"cb",
    x"27",
    x"82",
    x"ee",
    x"5f",
    x"89",
    x"0f",
    x"86",
    x"40",
    x"87",
    x"f1",
    x"88",
    x"02",
    x"58",
    x"c3",
    x"06",
    x"c5",
    x"4f",
    x"8a",
    x"cc",
    x"24",
    x"82",
    x"ee",
    x"5f",
    x"84",
    x"02",
    x"85",
    x"00",
    x"84",
    x"01",
    x"84",
    x"03",
    x"84",
    x"05",
    x"84",
    x"0e",
    x"1e",
    x"88",
    x"01",
    x"82",
    x"ee",
    x"5f",
    x"41",
    x"42",
    x"17",
    x"40",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"07",
    x"47",
    x"41",
    x"4c",
    x"41",
    x"47",
    x"41",
    x"21",
    x"00",
    x"e0",
    x"11",
    x"01",
    x"e0",
    x"01",
    x"fe",
    x"0f",
    x"36",
    x"00",
    x"ed",
    x"b0",
    x"31",
    x"00",
    x"e7",
    x"cd",
    x"38",
    x"01",
    x"e6",
    x"cf",
    x"4f",
    x"e6",
    x"0c",
    x"87",
    x"87",
    x"b1",
    x"cd",
    x"3b",
    x"01",
    x"cd",
    x"ad",
    x"59",
    x"3e",
    x"c3",
    x"21",
    x"4c",
    x"40",
    x"32",
    x"9a",
    x"fd",
    x"22",
    x"9b",
    x"fd",
    x"fb",
    x"01",
    x"01",
    x"e2",
    x"cd",
    x"47",
    x"00",
    x"18",
    x"fe",
    x"31",
    x"00",
    x"e7",
    x"cd",
    x"3e",
    x"01",
    x"01",
    x"01",
    x"c2",
    x"cd",
    x"47",
    x"00",
    x"2a",
    x"09",
    x"e0",
    x"23",
    x"22",
    x"09",
    x"e0",
    x"cb",
    x"45",
    x"28",
    x"18",
    x"21",
    x"80",
    x"e7",
    x"f9",
    x"3e",
    x"20",
    x"5e",
    x"2c",
    x"56",
    x"2c",
    x"4e",
    x"2c",
    x"46",
    x"2c",
    x"c5",
    x"d5",
    x"3d",
    x"20",
    x"f3",
    x"21",
    x"00",
    x"e7",
    x"18",
    x"03",
    x"21",
    x"80",
    x"e7",
    x"11",
    x"00",
    x"1b",
    x"01",
    x"80",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"21",
    x"61",
    x"e0",
    x"7e",
    x"11",
    x"00",
    x"01",
    x"d5",
    x"cd",
    x"af",
    x"41",
    x"3a",
    x"60",
    x"e0",
    x"86",
    x"77",
    x"d1",
    x"cd",
    x"b3",
    x"41",
    x"23",
    x"7e",
    x"11",
    x"20",
    x"01",
    x"d5",
    x"cd",
    x"af",
    x"41",
    x"3a",
    x"60",
    x"e0",
    x"cb",
    x"2f",
    x"86",
    x"77",
    x"d1",
    x"cd",
    x"b3",
    x"41",
    x"cd",
    x"20",
    x"90",
    x"3e",
    x"0f",
    x"1e",
    x"8f",
    x"cd",
    x"93",
    x"00",
    x"3e",
    x"0e",
    x"cd",
    x"96",
    x"00",
    x"32",
    x"30",
    x"e0",
    x"3e",
    x"0f",
    x"1e",
    x"cf",
    x"cd",
    x"93",
    x"00",
    x"3e",
    x"0e",
    x"cd",
    x"96",
    x"00",
    x"21",
    x"30",
    x"e0",
    x"a6",
    x"77",
    x"3e",
    x"08",
    x"cd",
    x"41",
    x"01",
    x"32",
    x"31",
    x"e0",
    x"07",
    x"cb",
    x"11",
    x"07",
    x"07",
    x"07",
    x"cb",
    x"11",
    x"3a",
    x"30",
    x"e0",
    x"1f",
    x"1f",
    x"a1",
    x"f6",
    x"fc",
    x"2f",
    x"32",
    x"20",
    x"e0",
    x"3e",
    x"05",
    x"cd",
    x"41",
    x"01",
    x"32",
    x"32",
    x"e0",
    x"f6",
    x"5f",
    x"4f",
    x"0f",
    x"a1",
    x"0f",
    x"4f",
    x"3a",
    x"30",
    x"e0",
    x"a1",
    x"4f",
    x"87",
    x"a1",
    x"07",
    x"07",
    x"07",
    x"4f",
    x"3a",
    x"31",
    x"e0",
    x"a1",
    x"f6",
    x"fe",
    x"2f",
    x"21",
    x"22",
    x"e0",
    x"4e",
    x"77",
    x"47",
    x"79",
    x"2f",
    x"a0",
    x"32",
    x"21",
    x"e0",
    x"3e",
    x"06",
    x"cd",
    x"41",
    x"01",
    x"e6",
    x"02",
    x"3e",
    x"ff",
    x"28",
    x"02",
    x"3e",
    x"9c",
    x"08",
    x"3e",
    x"07",
    x"cd",
    x"41",
    x"01",
    x"4f",
    x"2f",
    x"47",
    x"3a",
    x"24",
    x"e0",
    x"a0",
    x"47",
    x"08",
    x"a0",
    x"32",
    x"23",
    x"e0",
    x"79",
    x"f6",
    x"00",
    x"32",
    x"24",
    x"e0",
    x"21",
    x"0c",
    x"e0",
    x"3a",
    x"23",
    x"e0",
    x"e6",
    x"10",
    x"28",
    x"04",
    x"7e",
    x"ee",
    x"01",
    x"77",
    x"7e",
    x"3d",
    x"ca",
    x"5a",
    x"41",
    x"11",
    x"00",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"3a",
    x"00",
    x"e0",
    x"3d",
    x"cc",
    x"29",
    x"86",
    x"c3",
    x"44",
    x"40",
    x"21",
    x"00",
    x"00",
    x"39",
    x"eb",
    x"f9",
    x"e1",
    x"d5",
    x"f9",
    x"c9",
    x"21",
    x"00",
    x"00",
    x"39",
    x"5d",
    x"54",
    x"7d",
    x"e6",
    x"e0",
    x"6f",
    x"f9",
    x"e1",
    x"d5",
    x"f9",
    x"c9",
    x"21",
    x"00",
    x"e5",
    x"11",
    x"97",
    x"41",
    x"06",
    x"0b",
    x"7d",
    x"c6",
    x"1e",
    x"77",
    x"2c",
    x"74",
    x"6f",
    x"1a",
    x"77",
    x"2c",
    x"13",
    x"1a",
    x"77",
    x"23",
    x"13",
    x"10",
    x"ef",
    x"c9",
    x"d7",
    x"41",
    x"35",
    x"46",
    x"04",
    x"4d",
    x"03",
    x"80",
    x"5a",
    x"87",
    x"4e",
    x"53",
    x"0b",
    x"57",
    x"e3",
    x"48",
    x"93",
    x"81",
    x"5e",
    x"5e",
    x"48",
    x"58",
    x"00",
    x"00",
    x"0e",
    x"00",
    x"18",
    x"02",
    x"0e",
    x"20",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"eb",
    x"79",
    x"cd",
    x"4d",
    x"00",
    x"7c",
    x"c6",
    x"08",
    x"67",
    x"79",
    x"cd",
    x"4d",
    x"00",
    x"7c",
    x"c6",
    x"08",
    x"67",
    x"79",
    x"cd",
    x"4d",
    x"00",
    x"eb",
    x"c9",
    x"cd",
    x"f4",
    x"88",
    x"cd",
    x"6e",
    x"41",
    x"3a",
    x"21",
    x"e0",
    x"a7",
    x"20",
    x"02",
    x"18",
    x"f5",
    x"cd",
    x"a1",
    x"8a",
    x"3e",
    x"01",
    x"32",
    x"00",
    x"e0",
    x"32",
    x"50",
    x"e2",
    x"32",
    x"58",
    x"e2",
    x"32",
    x"60",
    x"e2",
    x"cd",
    x"1e",
    x"5a",
    x"cd",
    x"e1",
    x"88",
    x"21",
    x"f8",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"cd",
    x"6e",
    x"41",
    x"cd",
    x"e5",
    x"85",
    x"3a",
    x"50",
    x"e2",
    x"a7",
    x"20",
    x"f4",
    x"21",
    x"f8",
    x"45",
    x"cd",
    x"8f",
    x"8a",
    x"21",
    x"05",
    x"46",
    x"cd",
    x"7e",
    x"8a",
    x"06",
    x"5a",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"c1",
    x"10",
    x"f9",
    x"cd",
    x"41",
    x"81",
    x"21",
    x"05",
    x"46",
    x"cd",
    x"8f",
    x"8a",
    x"cd",
    x"f7",
    x"5a",
    x"cd",
    x"79",
    x"5a",
    x"21",
    x"74",
    x"e0",
    x"36",
    x"ff",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"60",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"20",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"a0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"c0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"3a",
    x"74",
    x"e0",
    x"a7",
    x"20",
    x"d3",
    x"3a",
    x"0d",
    x"e0",
    x"fe",
    x"03",
    x"ca",
    x"f2",
    x"43",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"20",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"20",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"e0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"a0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"c0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"00",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"cd",
    x"e5",
    x"85",
    x"3a",
    x"28",
    x"e0",
    x"fe",
    x"03",
    x"ca",
    x"ec",
    x"42",
    x"fe",
    x"0b",
    x"ca",
    x"ec",
    x"42",
    x"fe",
    x"09",
    x"ca",
    x"ec",
    x"42",
    x"21",
    x"17",
    x"e0",
    x"7e",
    x"a7",
    x"28",
    x"32",
    x"34",
    x"47",
    x"3d",
    x"20",
    x"09",
    x"21",
    x"0d",
    x"e0",
    x"7e",
    x"32",
    x"19",
    x"e0",
    x"36",
    x"00",
    x"78",
    x"fe",
    x"78",
    x"da",
    x"e4",
    x"42",
    x"3e",
    x"78",
    x"32",
    x"17",
    x"e0",
    x"3a",
    x"d7",
    x"e4",
    x"a7",
    x"ca",
    x"0c",
    x"43",
    x"c3",
    x"6c",
    x"42",
    x"3a",
    x"28",
    x"e0",
    x"d6",
    x"0b",
    x"c2",
    x"6c",
    x"42",
    x"af",
    x"32",
    x"17",
    x"e0",
    x"c3",
    x"6c",
    x"42",
    x"3a",
    x"10",
    x"e0",
    x"21",
    x"d7",
    x"e4",
    x"b6",
    x"21",
    x"92",
    x"e0",
    x"b6",
    x"c2",
    x"6c",
    x"42",
    x"3a",
    x"28",
    x"e0",
    x"fe",
    x"05",
    x"ca",
    x"6c",
    x"42",
    x"c3",
    x"2c",
    x"42",
    x"af",
    x"32",
    x"17",
    x"e0",
    x"32",
    x"18",
    x"e0",
    x"3a",
    x"19",
    x"e0",
    x"32",
    x"0d",
    x"e0",
    x"3a",
    x"0e",
    x"e0",
    x"a7",
    x"ca",
    x"47",
    x"43",
    x"21",
    x"05",
    x"46",
    x"cd",
    x"7e",
    x"8a",
    x"06",
    x"5a",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"20",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"c1",
    x"10",
    x"ed",
    x"cd",
    x"41",
    x"81",
    x"21",
    x"05",
    x"46",
    x"cd",
    x"8f",
    x"8a",
    x"c3",
    x"6c",
    x"42",
    x"21",
    x"0f",
    x"46",
    x"cd",
    x"7e",
    x"8a",
    x"06",
    x"f0",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"20",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"c1",
    x"10",
    x"f3",
    x"cd",
    x"e5",
    x"89",
    x"cd",
    x"03",
    x"8a",
    x"21",
    x"b3",
    x"45",
    x"06",
    x"04",
    x"c5",
    x"cd",
    x"7e",
    x"8a",
    x"c1",
    x"10",
    x"f9",
    x"cd",
    x"36",
    x"8b",
    x"21",
    x"51",
    x"19",
    x"11",
    x"f6",
    x"e0",
    x"01",
    x"05",
    x"03",
    x"cd",
    x"4f",
    x"8a",
    x"21",
    x"b1",
    x"19",
    x"11",
    x"f9",
    x"e0",
    x"01",
    x"05",
    x"03",
    x"cd",
    x"4f",
    x"8a",
    x"2a",
    x"f0",
    x"e0",
    x"7c",
    x"b5",
    x"28",
    x"0a",
    x"2a",
    x"f2",
    x"e0",
    x"7c",
    x"b5",
    x"28",
    x"53",
    x"cd",
    x"59",
    x"8b",
    x"21",
    x"13",
    x"1a",
    x"11",
    x"fe",
    x"e0",
    x"01",
    x"01",
    x"02",
    x"cd",
    x"4f",
    x"8a",
    x"21",
    x"15",
    x"1a",
    x"3e",
    x"8d",
    x"cd",
    x"4d",
    x"00",
    x"21",
    x"17",
    x"1a",
    x"3e",
    x"6b",
    x"cd",
    x"4d",
    x"00",
    x"3e",
    x"01",
    x"32",
    x"c0",
    x"e2",
    x"32",
    x"c8",
    x"e2",
    x"32",
    x"d0",
    x"e2",
    x"01",
    x"00",
    x"06",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"c1",
    x"3a",
    x"21",
    x"e0",
    x"a7",
    x"20",
    x"05",
    x"0b",
    x"79",
    x"b0",
    x"20",
    x"f0",
    x"af",
    x"32",
    x"c0",
    x"e2",
    x"32",
    x"c8",
    x"e2",
    x"32",
    x"d0",
    x"e2",
    x"32",
    x"00",
    x"e0",
    x"cd",
    x"6e",
    x"41",
    x"cd",
    x"e5",
    x"89",
    x"c3",
    x"d7",
    x"41",
    x"21",
    x"ef",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"18",
    x"c4",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"e0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"a0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"c0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"00",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"cd",
    x"e5",
    x"85",
    x"3a",
    x"0d",
    x"e0",
    x"a7",
    x"c2",
    x"f2",
    x"43",
    x"21",
    x"59",
    x"44",
    x"af",
    x"f5",
    x"e5",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"a0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"80",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"c0",
    x"e5",
    x"cd",
    x"64",
    x"41",
    x"11",
    x"40",
    x"e6",
    x"cd",
    x"64",
    x"41",
    x"cd",
    x"e5",
    x"85",
    x"e1",
    x"f1",
    x"be",
    x"3c",
    x"38",
    x"04",
    x"23",
    x"23",
    x"23",
    x"af",
    x"f5",
    x"e5",
    x"23",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"e9",
    x"96",
    x"a7",
    x"44",
    x"01",
    x"77",
    x"44",
    x"1e",
    x"a1",
    x"44",
    x"3c",
    x"aa",
    x"44",
    x"3c",
    x"b9",
    x"44",
    x"96",
    x"31",
    x"45",
    x"f0",
    x"fc",
    x"44",
    x"01",
    x"23",
    x"45",
    x"3c",
    x"a7",
    x"44",
    x"01",
    x"50",
    x"45",
    x"3a",
    x"a0",
    x"e0",
    x"fe",
    x"28",
    x"20",
    x"11",
    x"3e",
    x"01",
    x"32",
    x"88",
    x"e2",
    x"32",
    x"90",
    x"e2",
    x"32",
    x"98",
    x"e2",
    x"32",
    x"a3",
    x"e0",
    x"c3",
    x"29",
    x"44",
    x"3e",
    x"01",
    x"32",
    x"a0",
    x"e2",
    x"32",
    x"a8",
    x"e2",
    x"32",
    x"b8",
    x"e2",
    x"af",
    x"32",
    x"a3",
    x"e0",
    x"c3",
    x"29",
    x"44",
    x"21",
    x"6c",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"c3",
    x"29",
    x"44",
    x"21",
    x"13",
    x"19",
    x"11",
    x"a0",
    x"e0",
    x"01",
    x"01",
    x"01",
    x"cd",
    x"58",
    x"45",
    x"c3",
    x"29",
    x"44",
    x"3a",
    x"a3",
    x"e0",
    x"a7",
    x"21",
    x"8d",
    x"45",
    x"28",
    x"03",
    x"21",
    x"7d",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"21",
    x"a0",
    x"e0",
    x"7e",
    x"fe",
    x"28",
    x"20",
    x"02",
    x"36",
    x"64",
    x"cd",
    x"de",
    x"44",
    x"21",
    x"9b",
    x"45",
    x"cd",
    x"7e",
    x"8a",
    x"c3",
    x"29",
    x"44",
    x"11",
    x"a0",
    x"e0",
    x"1a",
    x"fe",
    x"64",
    x"30",
    x"10",
    x"21",
    x"88",
    x"19",
    x"af",
    x"cd",
    x"4d",
    x"00",
    x"21",
    x"89",
    x"19",
    x"01",
    x"02",
    x"01",
    x"c3",
    x"58",
    x"45",
    x"21",
    x"95",
    x"45",
    x"c3",
    x"7e",
    x"8a",
    x"3a",
    x"b8",
    x"e2",
    x"a7",
    x"20",
    x"2f",
    x"3a",
    x"b0",
    x"e2",
    x"a7",
    x"20",
    x"08",
    x"3a",
    x"a3",
    x"e0",
    x"ee",
    x"01",
    x"32",
    x"b0",
    x"e2",
    x"21",
    x"a0",
    x"e0",
    x"7e",
    x"a7",
    x"28",
    x"10",
    x"35",
    x"11",
    x"00",
    x"01",
    x"cd",
    x"a4",
    x"85",
    x"cd",
    x"de",
    x"44",
    x"18",
    x"0e",
    x"af",
    x"08",
    x"18",
    x"10",
    x"af",
    x"32",
    x"b0",
    x"e2",
    x"21",
    x"a4",
    x"45",
    x"cd",
    x"8f",
    x"8a",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"10",
    x"08",
    x"3a",
    x"a3",
    x"e0",
    x"a7",
    x"ca",
    x"29",
    x"44",
    x"21",
    x"a7",
    x"45",
    x"08",
    x"20",
    x"06",
    x"cd",
    x"7e",
    x"8a",
    x"c3",
    x"29",
    x"44",
    x"cd",
    x"8f",
    x"8a",
    x"c3",
    x"29",
    x"44",
    x"cd",
    x"03",
    x"8a",
    x"e1",
    x"e1",
    x"c3",
    x"2c",
    x"42",
    x"c5",
    x"1a",
    x"11",
    x"30",
    x"e0",
    x"a7",
    x"28",
    x"07",
    x"47",
    x"af",
    x"c6",
    x"01",
    x"27",
    x"10",
    x"fb",
    x"12",
    x"c1",
    x"c3",
    x"4f",
    x"8a",
    x"04",
    x"19",
    x"0e",
    x"7e",
    x"85",
    x"7d",
    x"72",
    x"75",
    x"82",
    x"27",
    x"7f",
    x"76",
    x"20",
    x"78",
    x"79",
    x"84",
    x"83",
    x"46",
    x"19",
    x"0d",
    x"13",
    x"10",
    x"05",
    x"03",
    x"09",
    x"01",
    x"0c",
    x"22",
    x"02",
    x"0f",
    x"0e",
    x"15",
    x"13",
    x"4a",
    x"19",
    x"05",
    x"72",
    x"7f",
    x"7e",
    x"85",
    x"83",
    x"88",
    x"19",
    x"03",
    x"61",
    x"60",
    x"60",
    x"8b",
    x"19",
    x"06",
    x"60",
    x"60",
    x"00",
    x"80",
    x"84",
    x"83",
    x"8b",
    x"19",
    x"02",
    x"a9",
    x"18",
    x"09",
    x"10",
    x"05",
    x"12",
    x"06",
    x"05",
    x"03",
    x"14",
    x"27",
    x"1e",
    x"e8",
    x"18",
    x"09",
    x"1c",
    x"12",
    x"05",
    x"13",
    x"15",
    x"0c",
    x"14",
    x"13",
    x"1c",
    x"43",
    x"19",
    x"0b",
    x"83",
    x"78",
    x"7f",
    x"84",
    x"83",
    x"00",
    x"76",
    x"79",
    x"82",
    x"75",
    x"74",
    x"a3",
    x"19",
    x"0e",
    x"7e",
    x"85",
    x"7d",
    x"72",
    x"75",
    x"82",
    x"00",
    x"7f",
    x"76",
    x"00",
    x"78",
    x"79",
    x"84",
    x"83",
    x"03",
    x"1a",
    x"0e",
    x"78",
    x"79",
    x"84",
    x"8b",
    x"7d",
    x"79",
    x"83",
    x"83",
    x"00",
    x"82",
    x"71",
    x"84",
    x"79",
    x"7f",
    x"12",
    x"1a",
    x"06",
    x"61",
    x"60",
    x"60",
    x"8d",
    x"60",
    x"6b",
    x"68",
    x"19",
    x"0a",
    x"77",
    x"71",
    x"7d",
    x"75",
    x"00",
    x"83",
    x"84",
    x"71",
    x"82",
    x"84",
    x"a9",
    x"19",
    x"07",
    x"12",
    x"05",
    x"01",
    x"04",
    x"19",
    x"25",
    x"1e",
    x"a8",
    x"19",
    x"09",
    x"77",
    x"71",
    x"7d",
    x"75",
    x"00",
    x"7f",
    x"86",
    x"75",
    x"82",
    x"19",
    x"18",
    x"04",
    x"08",
    x"09",
    x"07",
    x"08",
    x"3a",
    x"18",
    x"05",
    x"13",
    x"03",
    x"0f",
    x"12",
    x"05",
    x"99",
    x"18",
    x"05",
    x"13",
    x"03",
    x"0f",
    x"12",
    x"05",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"d0",
    x"e8",
    x"06",
    x"0d",
    x"cd",
    x"e1",
    x"8a",
    x"21",
    x"51",
    x"e0",
    x"7e",
    x"3c",
    x"fe",
    x"09",
    x"38",
    x"0c",
    x"11",
    x"52",
    x"e0",
    x"1a",
    x"3c",
    x"fe",
    x"10",
    x"38",
    x"01",
    x"af",
    x"12",
    x"af",
    x"77",
    x"3d",
    x"fa",
    x"1e",
    x"47",
    x"87",
    x"87",
    x"87",
    x"21",
    x"78",
    x"48",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"e5",
    x"dd",
    x"e1",
    x"6e",
    x"26",
    x"ef",
    x"11",
    x"d0",
    x"e8",
    x"01",
    x"0c",
    x"00",
    x"ed",
    x"b0",
    x"0e",
    x"14",
    x"09",
    x"0e",
    x"0c",
    x"ed",
    x"b0",
    x"dd",
    x"7e",
    x"01",
    x"06",
    x"0c",
    x"12",
    x"1c",
    x"3c",
    x"3c",
    x"10",
    x"fa",
    x"06",
    x"0c",
    x"d6",
    x"17",
    x"12",
    x"1c",
    x"3c",
    x"3c",
    x"10",
    x"fa",
    x"3a",
    x"51",
    x"e0",
    x"3d",
    x"e6",
    x"06",
    x"21",
    x"89",
    x"e3",
    x"85",
    x"6f",
    x"4e",
    x"2c",
    x"46",
    x"ed",
    x"43",
    x"87",
    x"e3",
    x"79",
    x"ed",
    x"44",
    x"dd",
    x"86",
    x"07",
    x"4f",
    x"dd",
    x"7e",
    x"02",
    x"c6",
    x"5a",
    x"6f",
    x"26",
    x"e3",
    x"06",
    x"05",
    x"71",
    x"2c",
    x"10",
    x"fc",
    x"dd",
    x"6e",
    x"02",
    x"26",
    x"e3",
    x"7d",
    x"fe",
    x"19",
    x"08",
    x"3a",
    x"52",
    x"e0",
    x"4f",
    x"e6",
    x"07",
    x"cb",
    x"45",
    x"28",
    x"0f",
    x"11",
    x"c0",
    x"48",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"79",
    x"fe",
    x"08",
    x"38",
    x"0f",
    x"18",
    x"2b",
    x"11",
    x"c8",
    x"48",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"79",
    x"fe",
    x"08",
    x"38",
    x"1e",
    x"1a",
    x"eb",
    x"21",
    x"2d",
    x"00",
    x"19",
    x"07",
    x"4f",
    x"06",
    x"05",
    x"cb",
    x"01",
    x"30",
    x"02",
    x"35",
    x"35",
    x"1a",
    x"a7",
    x"28",
    x"03",
    x"cd",
    x"c8",
    x"47",
    x"13",
    x"23",
    x"10",
    x"ef",
    x"c3",
    x"41",
    x"48",
    x"1a",
    x"eb",
    x"21",
    x"2d",
    x"00",
    x"19",
    x"07",
    x"4f",
    x"06",
    x"05",
    x"cb",
    x"01",
    x"30",
    x"02",
    x"34",
    x"34",
    x"1a",
    x"a7",
    x"28",
    x"03",
    x"cd",
    x"c8",
    x"47",
    x"13",
    x"23",
    x"10",
    x"ef",
    x"c3",
    x"41",
    x"48",
    x"3a",
    x"53",
    x"e0",
    x"3c",
    x"32",
    x"53",
    x"e0",
    x"11",
    x"00",
    x"e3",
    x"21",
    x"49",
    x"18",
    x"06",
    x"04",
    x"c5",
    x"1a",
    x"13",
    x"d5",
    x"e5",
    x"3d",
    x"28",
    x"6b",
    x"3d",
    x"28",
    x"57",
    x"18",
    x"39",
    x"e1",
    x"d1",
    x"23",
    x"23",
    x"c1",
    x"10",
    x"ec",
    x"3a",
    x"52",
    x"e0",
    x"11",
    x"ff",
    x"ff",
    x"cb",
    x"5f",
    x"28",
    x"04",
    x"11",
    x"01",
    x"00",
    x"2f",
    x"e6",
    x"07",
    x"21",
    x"b8",
    x"48",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"4e",
    x"cb",
    x"41",
    x"28",
    x"07",
    x"2a",
    x"8f",
    x"e3",
    x"19",
    x"22",
    x"8f",
    x"e3",
    x"cb",
    x"49",
    x"28",
    x"07",
    x"2a",
    x"8d",
    x"e3",
    x"19",
    x"22",
    x"8d",
    x"e3",
    x"c3",
    x"32",
    x"46",
    x"e5",
    x"01",
    x"02",
    x"00",
    x"eb",
    x"6b",
    x"26",
    x"ef",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"11",
    x"20",
    x"00",
    x"19",
    x"eb",
    x"6b",
    x"26",
    x"ef",
    x"01",
    x"02",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"18",
    x"ab",
    x"eb",
    x"21",
    x"d0",
    x"48",
    x"3a",
    x"53",
    x"e0",
    x"e6",
    x"04",
    x"28",
    x"15",
    x"23",
    x"23",
    x"23",
    x"23",
    x"18",
    x"0f",
    x"eb",
    x"21",
    x"d8",
    x"48",
    x"3a",
    x"53",
    x"e0",
    x"e6",
    x"04",
    x"28",
    x"04",
    x"23",
    x"23",
    x"23",
    x"23",
    x"e5",
    x"d5",
    x"01",
    x"02",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"eb",
    x"e1",
    x"23",
    x"23",
    x"0e",
    x"02",
    x"cd",
    x"5c",
    x"00",
    x"c3",
    x"3a",
    x"47",
    x"7e",
    x"d9",
    x"d6",
    x"08",
    x"fe",
    x"60",
    x"38",
    x"02",
    x"d6",
    x"60",
    x"47",
    x"c5",
    x"06",
    x"00",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"4f",
    x"21",
    x"d0",
    x"e8",
    x"09",
    x"eb",
    x"21",
    x"18",
    x"00",
    x"19",
    x"0e",
    x"03",
    x"ed",
    x"b0",
    x"0e",
    x"09",
    x"eb",
    x"09",
    x"eb",
    x"09",
    x"0e",
    x"03",
    x"ed",
    x"b0",
    x"08",
    x"30",
    x"06",
    x"08",
    x"21",
    x"00",
    x"e9",
    x"18",
    x"04",
    x"08",
    x"21",
    x"00",
    x"ec",
    x"3a",
    x"52",
    x"e0",
    x"e6",
    x"02",
    x"20",
    x"04",
    x"01",
    x"80",
    x"01",
    x"09",
    x"ed",
    x"4b",
    x"87",
    x"e3",
    x"09",
    x"eb",
    x"c1",
    x"78",
    x"e6",
    x"07",
    x"4f",
    x"87",
    x"81",
    x"87",
    x"87",
    x"87",
    x"87",
    x"30",
    x"01",
    x"14",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"21",
    x"00",
    x"e8",
    x"78",
    x"e6",
    x"f8",
    x"87",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"06",
    x"10",
    x"1a",
    x"13",
    x"b6",
    x"77",
    x"23",
    x"10",
    x"f9",
    x"0e",
    x"20",
    x"eb",
    x"ed",
    x"b0",
    x"d9",
    x"c9",
    x"dd",
    x"e5",
    x"cd",
    x"6e",
    x"41",
    x"dd",
    x"e1",
    x"dd",
    x"5e",
    x"03",
    x"dd",
    x"56",
    x"04",
    x"21",
    x"00",
    x"e8",
    x"01",
    x"c0",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"dd",
    x"5e",
    x"05",
    x"dd",
    x"56",
    x"06",
    x"21",
    x"d0",
    x"e8",
    x"01",
    x"0c",
    x"00",
    x"e5",
    x"d5",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"eb",
    x"e1",
    x"0e",
    x"0c",
    x"09",
    x"cd",
    x"5c",
    x"00",
    x"c3",
    x"32",
    x"46",
    x"81",
    x"a0",
    x"05",
    x"00",
    x"05",
    x"81",
    x"18",
    x"1f",
    x"8d",
    x"b8",
    x"0a",
    x"c0",
    x"05",
    x"8d",
    x"18",
    x"1f",
    x"c1",
    x"d0",
    x"0f",
    x"80",
    x"06",
    x"c1",
    x"18",
    x"2f",
    x"cd",
    x"e8",
    x"14",
    x"40",
    x"07",
    x"cd",
    x"18",
    x"2f",
    x"01",
    x"a0",
    x"19",
    x"00",
    x"0d",
    x"01",
    x"19",
    x"3f",
    x"0d",
    x"b8",
    x"1e",
    x"c0",
    x"0d",
    x"0d",
    x"19",
    x"3f",
    x"41",
    x"d0",
    x"23",
    x"80",
    x"0e",
    x"41",
    x"19",
    x"4f",
    x"4d",
    x"e8",
    x"28",
    x"40",
    x"0f",
    x"4d",
    x"19",
    x"4f",
    x"00",
    x"01",
    x"03",
    x"01",
    x"03",
    x"00",
    x"03",
    x"01",
    x"70",
    x"60",
    x"58",
    x"60",
    x"74",
    x"48",
    x"70",
    x"60",
    x"1c",
    x"0c",
    x"34",
    x"0c",
    x"5c",
    x"24",
    x"1c",
    x"0c",
    x"90",
    x"92",
    x"91",
    x"93",
    x"94",
    x"96",
    x"95",
    x"97",
    x"98",
    x"9a",
    x"99",
    x"9b",
    x"9c",
    x"9e",
    x"9d",
    x"9f",
    x"cd",
    x"6e",
    x"41",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"20",
    x"f7",
    x"3a",
    x"0d",
    x"e0",
    x"e6",
    x"01",
    x"c2",
    x"70",
    x"4b",
    x"21",
    x"96",
    x"e0",
    x"7e",
    x"3d",
    x"c2",
    x"48",
    x"49",
    x"3a",
    x"10",
    x"e0",
    x"d6",
    x"05",
    x"fe",
    x"06",
    x"d2",
    x"48",
    x"49",
    x"34",
    x"21",
    x"2c",
    x"e3",
    x"06",
    x"28",
    x"7e",
    x"a7",
    x"20",
    x"0a",
    x"2d",
    x"10",
    x"f9",
    x"3c",
    x"32",
    x"96",
    x"e0",
    x"c3",
    x"48",
    x"49",
    x"3e",
    x"01",
    x"32",
    x"00",
    x"e2",
    x"45",
    x"36",
    x"00",
    x"0e",
    x"03",
    x"78",
    x"d6",
    x"05",
    x"38",
    x"03",
    x"0c",
    x"18",
    x"f9",
    x"cd",
    x"b0",
    x"4a",
    x"46",
    x"7d",
    x"e6",
    x"3c",
    x"87",
    x"87",
    x"6f",
    x"26",
    x"e4",
    x"36",
    x"05",
    x"2c",
    x"2c",
    x"ed",
    x"5b",
    x"98",
    x"e0",
    x"73",
    x"2c",
    x"72",
    x"7d",
    x"c6",
    x"08",
    x"6f",
    x"36",
    x"00",
    x"2c",
    x"70",
    x"3a",
    x"14",
    x"e0",
    x"a7",
    x"ca",
    x"01",
    x"4a",
    x"3a",
    x"8c",
    x"e0",
    x"a7",
    x"c2",
    x"01",
    x"4a",
    x"21",
    x"d7",
    x"e4",
    x"3a",
    x"8a",
    x"e0",
    x"3d",
    x"be",
    x"da",
    x"01",
    x"4a",
    x"21",
    x"8e",
    x"e0",
    x"34",
    x"3a",
    x"82",
    x"e0",
    x"3d",
    x"be",
    x"d2",
    x"01",
    x"4a",
    x"36",
    x"00",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"03",
    x"26",
    x"e3",
    x"6f",
    x"7e",
    x"a7",
    x"20",
    x"09",
    x"2d",
    x"f2",
    x"77",
    x"49",
    x"2e",
    x"03",
    x"c3",
    x"77",
    x"49",
    x"f5",
    x"e5",
    x"21",
    x"91",
    x"e0",
    x"7e",
    x"34",
    x"e1",
    x"4d",
    x"e6",
    x"01",
    x"47",
    x"3a",
    x"28",
    x"e0",
    x"a7",
    x"28",
    x"02",
    x"06",
    x"00",
    x"c5",
    x"78",
    x"87",
    x"45",
    x"21",
    x"13",
    x"4b",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"eb",
    x"78",
    x"a7",
    x"28",
    x"09",
    x"fe",
    x"03",
    x"28",
    x"03",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"01",
    x"4f",
    x"c6",
    x"04",
    x"08",
    x"d5",
    x"cd",
    x"b0",
    x"4a",
    x"7d",
    x"e6",
    x"3c",
    x"87",
    x"87",
    x"c6",
    x"0c",
    x"32",
    x"30",
    x"e0",
    x"d1",
    x"c1",
    x"f1",
    x"3d",
    x"28",
    x"02",
    x"36",
    x"04",
    x"05",
    x"ca",
    x"01",
    x"4a",
    x"79",
    x"c6",
    x"07",
    x"6f",
    x"26",
    x"e3",
    x"06",
    x"03",
    x"0e",
    x"02",
    x"7e",
    x"a7",
    x"28",
    x"10",
    x"c5",
    x"d5",
    x"e5",
    x"45",
    x"08",
    x"4f",
    x"08",
    x"cd",
    x"b0",
    x"4a",
    x"e1",
    x"d1",
    x"c1",
    x"0d",
    x"28",
    x"03",
    x"2c",
    x"10",
    x"e9",
    x"3a",
    x"30",
    x"e0",
    x"6f",
    x"26",
    x"e4",
    x"79",
    x"ed",
    x"44",
    x"c6",
    x"02",
    x"77",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"01",
    x"ca",
    x"46",
    x"4a",
    x"3a",
    x"15",
    x"e0",
    x"a7",
    x"ca",
    x"e0",
    x"48",
    x"21",
    x"8f",
    x"e0",
    x"34",
    x"3a",
    x"88",
    x"e0",
    x"be",
    x"d2",
    x"e0",
    x"48",
    x"36",
    x"00",
    x"cd",
    x"c2",
    x"8a",
    x"26",
    x"e3",
    x"e6",
    x"02",
    x"28",
    x"10",
    x"2e",
    x"0f",
    x"7e",
    x"a7",
    x"20",
    x"13",
    x"2c",
    x"7d",
    x"fe",
    x"19",
    x"38",
    x"f6",
    x"2e",
    x"05",
    x"18",
    x"f2",
    x"2e",
    x"18",
    x"7e",
    x"a7",
    x"20",
    x"03",
    x"2d",
    x"18",
    x"f9",
    x"45",
    x"cd",
    x"90",
    x"4a",
    x"c3",
    x"e0",
    x"48",
    x"3a",
    x"16",
    x"e0",
    x"a7",
    x"ca",
    x"e0",
    x"48",
    x"21",
    x"90",
    x"e0",
    x"34",
    x"3a",
    x"86",
    x"e0",
    x"be",
    x"d2",
    x"e0",
    x"48",
    x"36",
    x"00",
    x"cd",
    x"c2",
    x"8a",
    x"26",
    x"e3",
    x"cb",
    x"4f",
    x"28",
    x"04",
    x"2e",
    x"19",
    x"18",
    x"02",
    x"2e",
    x"23",
    x"e6",
    x"80",
    x"28",
    x"12",
    x"7e",
    x"a7",
    x"20",
    x"18",
    x"2c",
    x"7d",
    x"fe",
    x"2d",
    x"38",
    x"f6",
    x"2e",
    x"19",
    x"18",
    x"f2",
    x"7e",
    x"a7",
    x"20",
    x"0a",
    x"2d",
    x"7d",
    x"fe",
    x"19",
    x"30",
    x"f6",
    x"2e",
    x"2c",
    x"18",
    x"f2",
    x"45",
    x"cd",
    x"90",
    x"4a",
    x"c3",
    x"e0",
    x"48",
    x"0e",
    x"03",
    x"78",
    x"d6",
    x"05",
    x"38",
    x"03",
    x"0c",
    x"18",
    x"f9",
    x"79",
    x"fe",
    x"08",
    x"30",
    x"05",
    x"11",
    x"ec",
    x"8b",
    x"18",
    x"03",
    x"11",
    x"c8",
    x"8b",
    x"21",
    x"d7",
    x"e4",
    x"3a",
    x"8a",
    x"e0",
    x"3d",
    x"be",
    x"d8",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"21",
    x"00",
    x"e4",
    x"7e",
    x"a7",
    x"ca",
    x"c2",
    x"4a",
    x"7d",
    x"c6",
    x"10",
    x"6f",
    x"18",
    x"f5",
    x"af",
    x"cb",
    x"39",
    x"1f",
    x"cb",
    x"39",
    x"0c",
    x"0c",
    x"71",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"73",
    x"2c",
    x"72",
    x"2c",
    x"77",
    x"2c",
    x"2c",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"2c",
    x"70",
    x"2c",
    x"77",
    x"2c",
    x"3a",
    x"93",
    x"e0",
    x"77",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"36",
    x"00",
    x"11",
    x"12",
    x"e0",
    x"79",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"3d",
    x"12",
    x"7d",
    x"21",
    x"82",
    x"e7",
    x"e6",
    x"f0",
    x"0f",
    x"0f",
    x"85",
    x"6f",
    x"0d",
    x"79",
    x"0f",
    x"0f",
    x"0f",
    x"77",
    x"2c",
    x"11",
    x"58",
    x"e0",
    x"79",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"77",
    x"c9",
    x"2e",
    x"8c",
    x"18",
    x"8c",
    x"af",
    x"32",
    x"0d",
    x"e0",
    x"3e",
    x"03",
    x"32",
    x"a9",
    x"e0",
    x"c3",
    x"e0",
    x"48",
    x"3a",
    x"d7",
    x"e4",
    x"a7",
    x"c2",
    x"e0",
    x"48",
    x"23",
    x"7e",
    x"fe",
    x"fe",
    x"28",
    x"e7",
    x"fe",
    x"fc",
    x"28",
    x"0a",
    x"2a",
    x"d0",
    x"e4",
    x"11",
    x"06",
    x"00",
    x"19",
    x"22",
    x"d0",
    x"e4",
    x"21",
    x"00",
    x"e4",
    x"22",
    x"d2",
    x"e4",
    x"e6",
    x"01",
    x"47",
    x"3a",
    x"d5",
    x"e4",
    x"11",
    x"ae",
    x"4c",
    x"87",
    x"80",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"32",
    x"d6",
    x"e4",
    x"11",
    x"d8",
    x"e4",
    x"2a",
    x"d0",
    x"e4",
    x"7e",
    x"12",
    x"23",
    x"13",
    x"7e",
    x"12",
    x"23",
    x"22",
    x"d0",
    x"e4",
    x"d9",
    x"34",
    x"34",
    x"3e",
    x"08",
    x"32",
    x"a9",
    x"e0",
    x"21",
    x"d4",
    x"e4",
    x"7e",
    x"d9",
    x"47",
    x"2a",
    x"9e",
    x"e0",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"fe",
    x"ff",
    x"28",
    x"a0",
    x"4f",
    x"78",
    x"e6",
    x"01",
    x"11",
    x"d8",
    x"e4",
    x"83",
    x"5f",
    x"1a",
    x"47",
    x"11",
    x"dc",
    x"e4",
    x"1a",
    x"b8",
    x"30",
    x"05",
    x"3c",
    x"12",
    x"c3",
    x"e0",
    x"48",
    x"af",
    x"12",
    x"d9",
    x"34",
    x"d9",
    x"7e",
    x"47",
    x"23",
    x"fe",
    x"e8",
    x"30",
    x"15",
    x"fe",
    x"e0",
    x"38",
    x"2a",
    x"11",
    x"d6",
    x"e4",
    x"1a",
    x"3d",
    x"fa",
    x"9c",
    x"4b",
    x"12",
    x"78",
    x"e6",
    x"03",
    x"4f",
    x"06",
    x"ff",
    x"18",
    x"23",
    x"11",
    x"a8",
    x"e0",
    x"1a",
    x"3d",
    x"c2",
    x"70",
    x"4b",
    x"12",
    x"3c",
    x"32",
    x"a5",
    x"e0",
    x"21",
    x"c0",
    x"e4",
    x"22",
    x"d2",
    x"e4",
    x"0e",
    x"ff",
    x"06",
    x"04",
    x"18",
    x"0a",
    x"78",
    x"07",
    x"07",
    x"e6",
    x"03",
    x"4f",
    x"78",
    x"e6",
    x"3f",
    x"47",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"2a",
    x"d2",
    x"e4",
    x"79",
    x"3c",
    x"3c",
    x"77",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"ed",
    x"5b",
    x"d0",
    x"e4",
    x"3a",
    x"d4",
    x"e4",
    x"1f",
    x"30",
    x"03",
    x"13",
    x"13",
    x"13",
    x"1a",
    x"13",
    x"77",
    x"2c",
    x"1a",
    x"13",
    x"77",
    x"2c",
    x"1a",
    x"77",
    x"2c",
    x"2c",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"2c",
    x"70",
    x"2c",
    x"77",
    x"2c",
    x"36",
    x"01",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"36",
    x"00",
    x"2c",
    x"2c",
    x"2c",
    x"22",
    x"d2",
    x"e4",
    x"7d",
    x"0f",
    x"0f",
    x"3d",
    x"21",
    x"80",
    x"e7",
    x"85",
    x"6f",
    x"11",
    x"58",
    x"e0",
    x"79",
    x"3c",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"77",
    x"c3",
    x"70",
    x"4b",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"b0",
    x"5f",
    x"80",
    x"b0",
    x"5f",
    x"00",
    x"08",
    x"00",
    x"b0",
    x"5f",
    x"80",
    x"b0",
    x"5f",
    x"00",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"08",
    x"b0",
    x"5f",
    x"00",
    x"b0",
    x"5f",
    x"00",
    x"08",
    x"08",
    x"b0",
    x"5f",
    x"80",
    x"b0",
    x"5f",
    x"80",
    x"08",
    x"08",
    x"c7",
    x"5f",
    x"80",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"08",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"9c",
    x"5f",
    x"00",
    x"b0",
    x"5f",
    x"00",
    x"08",
    x"00",
    x"9c",
    x"5f",
    x"80",
    x"b0",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"c7",
    x"5f",
    x"80",
    x"db",
    x"5f",
    x"80",
    x"08",
    x"00",
    x"db",
    x"5f",
    x"00",
    x"c7",
    x"5f",
    x"00",
    x"00",
    x"00",
    x"02",
    x"00",
    x"02",
    x"02",
    x"04",
    x"02",
    x"04",
    x"04",
    x"ff",
    x"fc",
    x"9d",
    x"49",
    x"9e",
    x"4a",
    x"e2",
    x"e1",
    x"a7",
    x"53",
    x"e2",
    x"e1",
    x"a8",
    x"54",
    x"ff",
    x"f1",
    x"00",
    x"48",
    x"e0",
    x"e1",
    x"01",
    x"4b",
    x"02",
    x"52",
    x"e0",
    x"e1",
    x"03",
    x"55",
    x"ff",
    x"f1",
    x"47",
    x"4c",
    x"e1",
    x"e1",
    x"46",
    x"4d",
    x"51",
    x"56",
    x"e1",
    x"e1",
    x"50",
    x"57",
    x"ff",
    x"f0",
    x"e2",
    x"e2",
    x"9c",
    x"9f",
    x"9b",
    x"a0",
    x"e2",
    x"e2",
    x"a6",
    x"a9",
    x"a5",
    x"aa",
    x"ff",
    x"f0",
    x"9a",
    x"a1",
    x"99",
    x"a2",
    x"a4",
    x"ab",
    x"e2",
    x"e2",
    x"e2",
    x"e2",
    x"a3",
    x"ac",
    x"e8",
    x"ff",
    x"fe",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"00",
    x"e4",
    x"dd",
    x"21",
    x"80",
    x"e7",
    x"06",
    x"0c",
    x"3a",
    x"a5",
    x"e0",
    x"a7",
    x"28",
    x"01",
    x"04",
    x"c5",
    x"e5",
    x"cd",
    x"28",
    x"4d",
    x"01",
    x"04",
    x"00",
    x"dd",
    x"09",
    x"e1",
    x"0e",
    x"10",
    x"09",
    x"c1",
    x"10",
    x"ef",
    x"c3",
    x"01",
    x"4d",
    x"e5",
    x"fd",
    x"e1",
    x"7e",
    x"a7",
    x"c8",
    x"3d",
    x"87",
    x"87",
    x"87",
    x"87",
    x"87",
    x"08",
    x"23",
    x"fd",
    x"7e",
    x"06",
    x"11",
    x"57",
    x"4d",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"47",
    x"7e",
    x"90",
    x"77",
    x"dc",
    x"5b",
    x"4d",
    x"23",
    x"23",
    x"23",
    x"7e",
    x"e6",
    x"7f",
    x"23",
    x"eb",
    x"21",
    x"12",
    x"4f",
    x"c3",
    x"f8",
    x"8a",
    x"04",
    x"07",
    x"0a",
    x"0e",
    x"23",
    x"5e",
    x"23",
    x"56",
    x"fd",
    x"35",
    x"0a",
    x"fa",
    x"66",
    x"4d",
    x"1b",
    x"1a",
    x"13",
    x"47",
    x"cb",
    x"7f",
    x"20",
    x"5b",
    x"23",
    x"4e",
    x"cb",
    x"09",
    x"cb",
    x"09",
    x"23",
    x"cb",
    x"77",
    x"20",
    x"1b",
    x"a9",
    x"cb",
    x"6f",
    x"7e",
    x"20",
    x"0a",
    x"3d",
    x"4f",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"0a",
    x"0d",
    x"18",
    x"07",
    x"3c",
    x"4f",
    x"e6",
    x"03",
    x"20",
    x"01",
    x"0c",
    x"79",
    x"e6",
    x"1f",
    x"77",
    x"2b",
    x"7e",
    x"e6",
    x"80",
    x"77",
    x"2b",
    x"72",
    x"2b",
    x"73",
    x"2b",
    x"78",
    x"e6",
    x"1f",
    x"87",
    x"87",
    x"86",
    x"77",
    x"f0",
    x"36",
    x"00",
    x"c9",
    x"e5",
    x"4d",
    x"ea",
    x"4d",
    x"ef",
    x"4d",
    x"fe",
    x"4d",
    x"06",
    x"4e",
    x"14",
    x"4e",
    x"32",
    x"4e",
    x"2b",
    x"4e",
    x"43",
    x"4e",
    x"4a",
    x"4e",
    x"63",
    x"4e",
    x"6d",
    x"4e",
    x"ad",
    x"4e",
    x"c1",
    x"4e",
    x"cf",
    x"4e",
    x"fb",
    x"4e",
    x"cb",
    x"77",
    x"20",
    x"09",
    x"e6",
    x"7f",
    x"e5",
    x"21",
    x"a8",
    x"4d",
    x"c3",
    x"f8",
    x"8a",
    x"e6",
    x"3f",
    x"fd",
    x"77",
    x"0a",
    x"18",
    x"8a",
    x"e1",
    x"72",
    x"2b",
    x"73",
    x"2b",
    x"c9",
    x"e1",
    x"18",
    x"81",
    x"fd",
    x"34",
    x"06",
    x"18",
    x"f8",
    x"fd",
    x"35",
    x"06",
    x"18",
    x"f3",
    x"1a",
    x"47",
    x"13",
    x"1a",
    x"13",
    x"fd",
    x"72",
    x"0f",
    x"fd",
    x"73",
    x"0e",
    x"57",
    x"58",
    x"18",
    x"e4",
    x"fd",
    x"56",
    x"0f",
    x"fd",
    x"5e",
    x"0e",
    x"18",
    x"dc",
    x"1a",
    x"13",
    x"47",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"b0",
    x"fd",
    x"77",
    x"04",
    x"18",
    x"c8",
    x"1a",
    x"47",
    x"13",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"20",
    x"05",
    x"fd",
    x"70",
    x"0d",
    x"18",
    x"bf",
    x"3e",
    x"1f",
    x"90",
    x"fd",
    x"77",
    x"0d",
    x"18",
    x"b7",
    x"1a",
    x"13",
    x"dd",
    x"77",
    x"00",
    x"18",
    x"b0",
    x"1a",
    x"13",
    x"fd",
    x"cb",
    x"04",
    x"7e",
    x"28",
    x"04",
    x"ed",
    x"44",
    x"c6",
    x"c0",
    x"dd",
    x"77",
    x"01",
    x"18",
    x"9f",
    x"1a",
    x"13",
    x"fd",
    x"77",
    x"06",
    x"18",
    x"98",
    x"1a",
    x"47",
    x"13",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"20",
    x"06",
    x"fd",
    x"70",
    x"05",
    x"c3",
    x"e2",
    x"4d",
    x"3e",
    x"1f",
    x"90",
    x"fd",
    x"77",
    x"05",
    x"c3",
    x"e2",
    x"4d",
    x"3a",
    x"dd",
    x"e4",
    x"a7",
    x"c2",
    x"e5",
    x"4d",
    x"c3",
    x"e2",
    x"4d",
    x"3a",
    x"93",
    x"e0",
    x"fd",
    x"77",
    x"0b",
    x"dd",
    x"e5",
    x"e1",
    x"7e",
    x"c6",
    x"30",
    x"77",
    x"3a",
    x"0d",
    x"e0",
    x"fe",
    x"02",
    x"20",
    x"1e",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"20",
    x"18",
    x"2c",
    x"7e",
    x"fd",
    x"cb",
    x"04",
    x"7e",
    x"28",
    x"04",
    x"ed",
    x"44",
    x"c6",
    x"c0",
    x"d6",
    x"70",
    x"f2",
    x"9a",
    x"4e",
    x"c6",
    x"50",
    x"c6",
    x"20",
    x"c3",
    x"34",
    x"4e",
    x"fd",
    x"7e",
    x"09",
    x"21",
    x"2d",
    x"e3",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"18",
    x"91",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"20",
    x"08",
    x"3a",
    x"0d",
    x"e0",
    x"fe",
    x"02",
    x"ca",
    x"e2",
    x"4d",
    x"11",
    x"ee",
    x"5f",
    x"c3",
    x"e2",
    x"4d",
    x"3a",
    x"85",
    x"e0",
    x"a7",
    x"ca",
    x"e2",
    x"4d",
    x"fd",
    x"36",
    x"06",
    x"02",
    x"c3",
    x"e2",
    x"4d",
    x"21",
    x"20",
    x"e1",
    x"7e",
    x"a7",
    x"c2",
    x"e2",
    x"4d",
    x"36",
    x"01",
    x"23",
    x"dd",
    x"7e",
    x"01",
    x"77",
    x"23",
    x"36",
    x"00",
    x"e1",
    x"e5",
    x"7d",
    x"e6",
    x"f0",
    x"32",
    x"25",
    x"e1",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"f6",
    x"09",
    x"fd",
    x"77",
    x"04",
    x"3e",
    x"01",
    x"32",
    x"b8",
    x"e1",
    x"c3",
    x"dc",
    x"4d",
    x"fd",
    x"7e",
    x"00",
    x"fe",
    x"02",
    x"ca",
    x"e2",
    x"4d",
    x"c3",
    x"fe",
    x"4d",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"c2",
    x"ef",
    x"4d",
    x"13",
    x"13",
    x"c3",
    x"e2",
    x"4d",
    x"34",
    x"4f",
    x"d9",
    x"4f",
    x"3f",
    x"50",
    x"c1",
    x"50",
    x"49",
    x"51",
    x"76",
    x"51",
    x"d5",
    x"4f",
    x"93",
    x"51",
    x"b6",
    x"51",
    x"94",
    x"52",
    x"83",
    x"51",
    x"ac",
    x"52",
    x"ce",
    x"51",
    x"fd",
    x"51",
    x"77",
    x"52",
    x"93",
    x"52",
    x"6e",
    x"51",
    x"eb",
    x"7e",
    x"47",
    x"23",
    x"7e",
    x"23",
    x"e6",
    x"03",
    x"28",
    x"5c",
    x"0f",
    x"0f",
    x"0f",
    x"80",
    x"11",
    x"80",
    x"9f",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"86",
    x"c6",
    x"08",
    x"47",
    x"fa",
    x"5a",
    x"4f",
    x"fe",
    x"10",
    x"38",
    x"10",
    x"e6",
    x"f0",
    x"18",
    x"02",
    x"f6",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"dd",
    x"86",
    x"00",
    x"dd",
    x"77",
    x"00",
    x"78",
    x"e6",
    x"0f",
    x"d6",
    x"08",
    x"77",
    x"23",
    x"7b",
    x"c6",
    x"08",
    x"e6",
    x"1f",
    x"47",
    x"7b",
    x"e6",
    x"e0",
    x"b0",
    x"5f",
    x"1a",
    x"86",
    x"c6",
    x"08",
    x"47",
    x"fa",
    x"88",
    x"4f",
    x"fe",
    x"10",
    x"38",
    x"10",
    x"e6",
    x"f0",
    x"18",
    x"02",
    x"f6",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"dd",
    x"86",
    x"01",
    x"dd",
    x"77",
    x"01",
    x"78",
    x"e6",
    x"0f",
    x"d6",
    x"08",
    x"77",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"7f",
    x"fe",
    x"02",
    x"28",
    x"0e",
    x"fd",
    x"7e",
    x"05",
    x"3c",
    x"3c",
    x"e6",
    x"1c",
    x"47",
    x"08",
    x"80",
    x"dd",
    x"77",
    x"02",
    x"c9",
    x"fd",
    x"7e",
    x"05",
    x"3c",
    x"3c",
    x"e6",
    x"1c",
    x"47",
    x"fd",
    x"be",
    x"0d",
    x"20",
    x"06",
    x"08",
    x"80",
    x"dd",
    x"77",
    x"02",
    x"c9",
    x"fd",
    x"7e",
    x"0d",
    x"e6",
    x"1c",
    x"b8",
    x"28",
    x"05",
    x"04",
    x"fd",
    x"70",
    x"0d",
    x"c9",
    x"fd",
    x"35",
    x"0d",
    x"c9",
    x"26",
    x"ff",
    x"18",
    x"02",
    x"26",
    x"00",
    x"fd",
    x"46",
    x"0d",
    x"78",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"05",
    x"78",
    x"3c",
    x"e6",
    x"1f",
    x"47",
    x"1a",
    x"4f",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"05",
    x"79",
    x"3c",
    x"e6",
    x"1f",
    x"4f",
    x"79",
    x"90",
    x"28",
    x"27",
    x"e6",
    x"1f",
    x"fe",
    x"10",
    x"30",
    x"0a",
    x"0d",
    x"79",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"0b",
    x"0d",
    x"18",
    x"08",
    x"0c",
    x"79",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"01",
    x"0c",
    x"79",
    x"e6",
    x"1f",
    x"12",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"24",
    x"ca",
    x"34",
    x"4f",
    x"c3",
    x"9a",
    x"4f",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"c9",
    x"06",
    x"04",
    x"11",
    x"ff",
    x"e2",
    x"13",
    x"1a",
    x"a7",
    x"20",
    x"02",
    x"10",
    x"f9",
    x"7b",
    x"32",
    x"a7",
    x"e0",
    x"87",
    x"87",
    x"87",
    x"87",
    x"c6",
    x"48",
    x"32",
    x"31",
    x"e3",
    x"c9",
    x"d5",
    x"fd",
    x"e5",
    x"e1",
    x"7e",
    x"3d",
    x"cc",
    x"25",
    x"50",
    x"fd",
    x"7e",
    x"09",
    x"fe",
    x"2d",
    x"30",
    x"52",
    x"c6",
    x"2d",
    x"6f",
    x"26",
    x"e3",
    x"5e",
    x"c6",
    x"2d",
    x"6f",
    x"56",
    x"dd",
    x"66",
    x"00",
    x"dd",
    x"6e",
    x"01",
    x"cd",
    x"d4",
    x"52",
    x"67",
    x"78",
    x"81",
    x"38",
    x"04",
    x"fe",
    x"08",
    x"38",
    x"2a",
    x"44",
    x"d1",
    x"1a",
    x"4f",
    x"90",
    x"28",
    x"18",
    x"e6",
    x"1f",
    x"fe",
    x"10",
    x"30",
    x"0a",
    x"0d",
    x"79",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"0b",
    x"0d",
    x"18",
    x"08",
    x"0c",
    x"79",
    x"2f",
    x"e6",
    x"03",
    x"20",
    x"01",
    x"0c",
    x"79",
    x"e6",
    x"1f",
    x"12",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"c3",
    x"34",
    x"4f",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"dd",
    x"72",
    x"00",
    x"dd",
    x"73",
    x"01",
    x"d1",
    x"c9",
    x"2c",
    x"36",
    x"00",
    x"11",
    x"b9",
    x"50",
    x"2c",
    x"73",
    x"2c",
    x"72",
    x"dd",
    x"56",
    x"00",
    x"dd",
    x"5e",
    x"01",
    x"cd",
    x"8a",
    x"59",
    x"fd",
    x"77",
    x"0d",
    x"d1",
    x"c9",
    x"88",
    x"02",
    x"84",
    x"06",
    x"cf",
    x"48",
    x"84",
    x"05",
    x"fd",
    x"7e",
    x"00",
    x"3d",
    x"28",
    x"46",
    x"fd",
    x"36",
    x"01",
    x"88",
    x"fd",
    x"34",
    x"04",
    x"13",
    x"13",
    x"af",
    x"12",
    x"26",
    x"e3",
    x"fd",
    x"7e",
    x"09",
    x"6f",
    x"fe",
    x"05",
    x"30",
    x"0b",
    x"dd",
    x"7e",
    x"03",
    x"fe",
    x"04",
    x"20",
    x"04",
    x"36",
    x"02",
    x"18",
    x"02",
    x"36",
    x"01",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"01",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"00",
    x"fd",
    x"7e",
    x"00",
    x"3d",
    x"3d",
    x"fe",
    x"03",
    x"28",
    x"3a",
    x"d0",
    x"21",
    x"14",
    x"e0",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"34",
    x"c9",
    x"fd",
    x"36",
    x"00",
    x"00",
    x"3e",
    x"05",
    x"32",
    x"28",
    x"e0",
    x"21",
    x"d7",
    x"e4",
    x"35",
    x"21",
    x"c0",
    x"e4",
    x"36",
    x"01",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"01",
    x"55",
    x"8c",
    x"71",
    x"2c",
    x"70",
    x"2c",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"80",
    x"77",
    x"7d",
    x"c6",
    x"06",
    x"6f",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"32",
    x"a5",
    x"e0",
    x"c9",
    x"fd",
    x"7e",
    x"09",
    x"21",
    x"15",
    x"e0",
    x"fe",
    x"19",
    x"38",
    x"01",
    x"23",
    x"34",
    x"c9",
    x"3a",
    x"51",
    x"e0",
    x"e6",
    x"01",
    x"c0",
    x"fd",
    x"7e",
    x"09",
    x"4f",
    x"26",
    x"e3",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"be",
    x"01",
    x"20",
    x"0b",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"be",
    x"00",
    x"20",
    x"01",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"c9",
    x"af",
    x"32",
    x"a5",
    x"e0",
    x"3c",
    x"32",
    x"a8",
    x"e0",
    x"21",
    x"d7",
    x"e4",
    x"35",
    x"fd",
    x"36",
    x"00",
    x"00",
    x"dd",
    x"36",
    x"00",
    x"e0",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"c0",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"f6",
    x"08",
    x"fd",
    x"77",
    x"04",
    x"18",
    x"07",
    x"fd",
    x"36",
    x"01",
    x"88",
    x"fd",
    x"34",
    x"04",
    x"fd",
    x"36",
    x"06",
    x"00",
    x"26",
    x"e3",
    x"fd",
    x"6e",
    x"09",
    x"36",
    x"00",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"01",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"00",
    x"c9",
    x"fd",
    x"7e",
    x"01",
    x"fe",
    x"09",
    x"d0",
    x"3e",
    x"01",
    x"32",
    x"08",
    x"e2",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"fd",
    x"77",
    x"04",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"f6",
    x"0d",
    x"fd",
    x"77",
    x"04",
    x"fd",
    x"36",
    x"06",
    x"00",
    x"26",
    x"e3",
    x"fd",
    x"7e",
    x"09",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"01",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"dd",
    x"77",
    x"00",
    x"3e",
    x"3c",
    x"32",
    x"97",
    x"e0",
    x"fd",
    x"7e",
    x"09",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"21",
    x"97",
    x"e0",
    x"35",
    x"28",
    x"11",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"10",
    x"fd",
    x"7e",
    x"0c",
    x"20",
    x"03",
    x"3a",
    x"5c",
    x"e0",
    x"dd",
    x"77",
    x"03",
    x"c9",
    x"af",
    x"fd",
    x"77",
    x"01",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"fd",
    x"77",
    x"04",
    x"3a",
    x"5c",
    x"e0",
    x"dd",
    x"77",
    x"03",
    x"dd",
    x"36",
    x"02",
    x"80",
    x"eb",
    x"7d",
    x"e6",
    x"f0",
    x"6f",
    x"e5",
    x"11",
    x"a0",
    x"e4",
    x"01",
    x"10",
    x"00",
    x"ed",
    x"b0",
    x"e1",
    x"7d",
    x"0e",
    x"10",
    x"ed",
    x"b0",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"c6",
    x"80",
    x"6f",
    x"26",
    x"e7",
    x"e5",
    x"11",
    x"a8",
    x"e7",
    x"0e",
    x"04",
    x"ed",
    x"b0",
    x"e1",
    x"0e",
    x"04",
    x"ed",
    x"b0",
    x"3e",
    x"ff",
    x"32",
    x"a9",
    x"e4",
    x"32",
    x"b9",
    x"e4",
    x"2a",
    x"9a",
    x"e0",
    x"22",
    x"a2",
    x"e4",
    x"2a",
    x"9c",
    x"e0",
    x"22",
    x"b2",
    x"e4",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"34",
    x"3e",
    x"01",
    x"32",
    x"08",
    x"e2",
    x"c9",
    x"eb",
    x"2d",
    x"2d",
    x"56",
    x"2d",
    x"5e",
    x"2d",
    x"1a",
    x"87",
    x"87",
    x"77",
    x"2c",
    x"1a",
    x"13",
    x"73",
    x"2c",
    x"72",
    x"2c",
    x"2c",
    x"eb",
    x"fd",
    x"34",
    x"04",
    x"fd",
    x"36",
    x"06",
    x"00",
    x"c9",
    x"c9",
    x"3a",
    x"20",
    x"e1",
    x"a7",
    x"28",
    x"05",
    x"fd",
    x"36",
    x"01",
    x"7f",
    x"c9",
    x"fd",
    x"36",
    x"01",
    x"00",
    x"fd",
    x"7e",
    x"04",
    x"e6",
    x"80",
    x"fd",
    x"77",
    x"04",
    x"c9",
    x"d5",
    x"eb",
    x"2d",
    x"2d",
    x"56",
    x"2d",
    x"5e",
    x"2d",
    x"36",
    x"7f",
    x"eb",
    x"dd",
    x"7e",
    x"00",
    x"96",
    x"f2",
    x"c0",
    x"52",
    x"ed",
    x"44",
    x"fe",
    x"04",
    x"d9",
    x"d1",
    x"d2",
    x"34",
    x"4f",
    x"d9",
    x"eb",
    x"36",
    x"00",
    x"2c",
    x"13",
    x"73",
    x"2c",
    x"72",
    x"d9",
    x"c3",
    x"34",
    x"4f",
    x"7c",
    x"c6",
    x"20",
    x"67",
    x"7a",
    x"c6",
    x"20",
    x"94",
    x"30",
    x"13",
    x"ed",
    x"44",
    x"4f",
    x"7b",
    x"95",
    x"30",
    x"07",
    x"ed",
    x"44",
    x"47",
    x"26",
    x"18",
    x"18",
    x"14",
    x"47",
    x"26",
    x"00",
    x"18",
    x"0f",
    x"4f",
    x"7b",
    x"95",
    x"30",
    x"07",
    x"ed",
    x"44",
    x"47",
    x"26",
    x"10",
    x"18",
    x"03",
    x"47",
    x"26",
    x"08",
    x"78",
    x"b9",
    x"38",
    x"06",
    x"41",
    x"4f",
    x"3e",
    x"04",
    x"84",
    x"67",
    x"79",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"6f",
    x"cb",
    x"3f",
    x"b8",
    x"30",
    x"0b",
    x"24",
    x"85",
    x"b8",
    x"30",
    x"06",
    x"24",
    x"87",
    x"b8",
    x"30",
    x"01",
    x"24",
    x"7c",
    x"21",
    x"2b",
    x"53",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"c9",
    x"00",
    x"01",
    x"02",
    x"04",
    x"08",
    x"06",
    x"05",
    x"04",
    x"10",
    x"0e",
    x"0d",
    x"0c",
    x"08",
    x"09",
    x"0a",
    x"0c",
    x"10",
    x"11",
    x"12",
    x"14",
    x"18",
    x"16",
    x"15",
    x"14",
    x"00",
    x"1e",
    x"1d",
    x"1c",
    x"18",
    x"19",
    x"1a",
    x"1c",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"57",
    x"53",
    x"3a",
    x"28",
    x"e0",
    x"c3",
    x"f8",
    x"8a",
    x"6f",
    x"53",
    x"ae",
    x"53",
    x"36",
    x"54",
    x"8e",
    x"55",
    x"34",
    x"56",
    x"80",
    x"56",
    x"6f",
    x"53",
    x"6f",
    x"53",
    x"04",
    x"54",
    x"58",
    x"55",
    x"03",
    x"55",
    x"e4",
    x"55",
    x"21",
    x"b4",
    x"e7",
    x"7e",
    x"fe",
    x"e0",
    x"28",
    x"d4",
    x"23",
    x"11",
    x"29",
    x"e0",
    x"3a",
    x"20",
    x"e0",
    x"a7",
    x"ca",
    x"4b",
    x"53",
    x"fe",
    x"03",
    x"ca",
    x"4b",
    x"53",
    x"0f",
    x"da",
    x"9c",
    x"53",
    x"7e",
    x"fe",
    x"b8",
    x"d2",
    x"4b",
    x"53",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"01",
    x"3c",
    x"86",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"7e",
    x"fe",
    x"08",
    x"da",
    x"4b",
    x"53",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"01",
    x"3d",
    x"3d",
    x"86",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"b5",
    x"e7",
    x"11",
    x"29",
    x"e0",
    x"3a",
    x"20",
    x"e0",
    x"a7",
    x"ca",
    x"4b",
    x"53",
    x"fe",
    x"03",
    x"ca",
    x"4b",
    x"53",
    x"0f",
    x"da",
    x"dc",
    x"53",
    x"7e",
    x"fe",
    x"aa",
    x"d2",
    x"4b",
    x"53",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"01",
    x"3c",
    x"86",
    x"77",
    x"2d",
    x"2d",
    x"2d",
    x"2d",
    x"c6",
    x"0d",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"7e",
    x"fe",
    x"08",
    x"da",
    x"4b",
    x"53",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"01",
    x"3d",
    x"3d",
    x"86",
    x"77",
    x"2d",
    x"2d",
    x"2d",
    x"2d",
    x"c6",
    x"0d",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"3e",
    x"08",
    x"32",
    x"28",
    x"e0",
    x"af",
    x"32",
    x"c0",
    x"e1",
    x"3a",
    x"63",
    x"e0",
    x"32",
    x"60",
    x"e0",
    x"21",
    x"b4",
    x"e7",
    x"34",
    x"7e",
    x"2c",
    x"2c",
    x"fe",
    x"a3",
    x"28",
    x"1b",
    x"11",
    x"29",
    x"e0",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"03",
    x"c2",
    x"4b",
    x"53",
    x"7e",
    x"a7",
    x"ca",
    x"4b",
    x"53",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"2c",
    x"36",
    x"0f",
    x"c3",
    x"4b",
    x"53",
    x"36",
    x"00",
    x"af",
    x"32",
    x"28",
    x"e0",
    x"32",
    x"18",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"c0",
    x"e1",
    x"7e",
    x"a7",
    x"20",
    x"01",
    x"34",
    x"af",
    x"32",
    x"b8",
    x"e1",
    x"3e",
    x"f0",
    x"32",
    x"60",
    x"e0",
    x"21",
    x"b4",
    x"e7",
    x"7e",
    x"fe",
    x"78",
    x"28",
    x"31",
    x"35",
    x"23",
    x"3a",
    x"21",
    x"e1",
    x"be",
    x"28",
    x"06",
    x"38",
    x"03",
    x"34",
    x"18",
    x"01",
    x"35",
    x"23",
    x"3a",
    x"25",
    x"e1",
    x"5f",
    x"16",
    x"e4",
    x"1a",
    x"a7",
    x"28",
    x"8d",
    x"11",
    x"29",
    x"e0",
    x"1a",
    x"3c",
    x"12",
    x"e6",
    x"03",
    x"20",
    x"06",
    x"7e",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"21",
    x"22",
    x"e1",
    x"36",
    x"00",
    x"c3",
    x"4b",
    x"53",
    x"2c",
    x"2c",
    x"7e",
    x"a7",
    x"20",
    x"d8",
    x"21",
    x"20",
    x"e1",
    x"36",
    x"03",
    x"7d",
    x"c6",
    x"05",
    x"6f",
    x"7e",
    x"11",
    x"a6",
    x"e0",
    x"12",
    x"13",
    x"26",
    x"e4",
    x"3c",
    x"6f",
    x"36",
    x"00",
    x"2c",
    x"01",
    x"f8",
    x"5f",
    x"71",
    x"2c",
    x"70",
    x"2c",
    x"36",
    x"00",
    x"7d",
    x"c6",
    x"05",
    x"6f",
    x"7e",
    x"12",
    x"21",
    x"b4",
    x"e7",
    x"11",
    x"b0",
    x"e7",
    x"01",
    x"03",
    x"00",
    x"ed",
    x"b0",
    x"3e",
    x"08",
    x"12",
    x"13",
    x"3e",
    x"e0",
    x"12",
    x"21",
    x"28",
    x"e0",
    x"36",
    x"0a",
    x"af",
    x"32",
    x"c0",
    x"e1",
    x"32",
    x"29",
    x"e0",
    x"3c",
    x"21",
    x"c0",
    x"e4",
    x"77",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"01",
    x"55",
    x"8c",
    x"71",
    x"2c",
    x"70",
    x"2c",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"80",
    x"77",
    x"7d",
    x"c6",
    x"06",
    x"6f",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"21",
    x"f0",
    x"54",
    x"cd",
    x"7e",
    x"8a",
    x"c3",
    x"4b",
    x"53",
    x"85",
    x"19",
    x"10",
    x"76",
    x"79",
    x"77",
    x"78",
    x"84",
    x"75",
    x"82",
    x"00",
    x"73",
    x"71",
    x"80",
    x"84",
    x"85",
    x"82",
    x"75",
    x"74",
    x"21",
    x"29",
    x"e0",
    x"34",
    x"7e",
    x"fe",
    x"78",
    x"30",
    x"1b",
    x"fe",
    x"1e",
    x"20",
    x"0b",
    x"3e",
    x"01",
    x"32",
    x"38",
    x"e2",
    x"32",
    x"40",
    x"e2",
    x"32",
    x"48",
    x"e2",
    x"3a",
    x"a6",
    x"e0",
    x"6f",
    x"2c",
    x"26",
    x"e4",
    x"36",
    x"7f",
    x"c3",
    x"4b",
    x"53",
    x"3a",
    x"a6",
    x"e0",
    x"6f",
    x"2c",
    x"26",
    x"e4",
    x"36",
    x"00",
    x"21",
    x"f0",
    x"54",
    x"cd",
    x"8f",
    x"8a",
    x"3e",
    x"04",
    x"32",
    x"28",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"3e",
    x"09",
    x"32",
    x"28",
    x"e0",
    x"3e",
    x"01",
    x"32",
    x"18",
    x"e0",
    x"32",
    x"d8",
    x"e1",
    x"32",
    x"28",
    x"e2",
    x"32",
    x"30",
    x"e2",
    x"21",
    x"a5",
    x"e0",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"21",
    x"a6",
    x"e0",
    x"34",
    x"7e",
    x"fe",
    x"3c",
    x"38",
    x"09",
    x"3a",
    x"d7",
    x"e4",
    x"21",
    x"92",
    x"e0",
    x"b6",
    x"28",
    x"17",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"03",
    x"c2",
    x"7b",
    x"55",
    x"21",
    x"b2",
    x"e7",
    x"7e",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"2c",
    x"36",
    x"0f",
    x"c3",
    x"6f",
    x"53",
    x"3a",
    x"b4",
    x"e7",
    x"fe",
    x"e0",
    x"ca",
    x"df",
    x"55",
    x"3e",
    x"03",
    x"32",
    x"28",
    x"e0",
    x"21",
    x"b2",
    x"e7",
    x"7e",
    x"a7",
    x"28",
    x"0f",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"03",
    x"20",
    x"24",
    x"7e",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"18",
    x"1c",
    x"2d",
    x"7e",
    x"fe",
    x"67",
    x"28",
    x"08",
    x"38",
    x"03",
    x"35",
    x"18",
    x"11",
    x"34",
    x"18",
    x"0e",
    x"3a",
    x"b5",
    x"e7",
    x"fe",
    x"5a",
    x"20",
    x"07",
    x"2d",
    x"7e",
    x"fe",
    x"a3",
    x"28",
    x"14",
    x"34",
    x"21",
    x"b5",
    x"e7",
    x"7e",
    x"fe",
    x"5a",
    x"ca",
    x"4b",
    x"53",
    x"38",
    x"04",
    x"35",
    x"c3",
    x"4b",
    x"53",
    x"34",
    x"c3",
    x"4b",
    x"53",
    x"3e",
    x"01",
    x"32",
    x"28",
    x"e0",
    x"af",
    x"32",
    x"18",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"3e",
    x"0b",
    x"32",
    x"28",
    x"e0",
    x"21",
    x"b2",
    x"e7",
    x"7e",
    x"a7",
    x"28",
    x"11",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"03",
    x"c2",
    x"4b",
    x"53",
    x"7e",
    x"c6",
    x"04",
    x"e6",
    x"1f",
    x"77",
    x"c3",
    x"4b",
    x"53",
    x"2d",
    x"7e",
    x"fe",
    x"60",
    x"28",
    x"0a",
    x"38",
    x"04",
    x"35",
    x"c3",
    x"4b",
    x"53",
    x"34",
    x"c3",
    x"4b",
    x"53",
    x"2d",
    x"7e",
    x"fe",
    x"a3",
    x"28",
    x"04",
    x"34",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"b0",
    x"e7",
    x"11",
    x"b4",
    x"e7",
    x"01",
    x"04",
    x"00",
    x"ed",
    x"b0",
    x"3e",
    x"e0",
    x"32",
    x"b0",
    x"e7",
    x"af",
    x"32",
    x"28",
    x"e0",
    x"32",
    x"17",
    x"e0",
    x"af",
    x"32",
    x"18",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"11",
    x"a7",
    x"e0",
    x"1a",
    x"6f",
    x"26",
    x"e3",
    x"7e",
    x"a7",
    x"c2",
    x"66",
    x"56",
    x"1b",
    x"1a",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"c6",
    x"80",
    x"6f",
    x"26",
    x"e7",
    x"11",
    x"b0",
    x"e7",
    x"7e",
    x"fe",
    x"68",
    x"f5",
    x"2c",
    x"c6",
    x"10",
    x"12",
    x"1c",
    x"7e",
    x"2c",
    x"12",
    x"f1",
    x"d2",
    x"4b",
    x"53",
    x"1c",
    x"7e",
    x"e6",
    x"1f",
    x"12",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"b0",
    x"e7",
    x"35",
    x"f2",
    x"4b",
    x"53",
    x"3e",
    x"01",
    x"32",
    x"17",
    x"e0",
    x"3e",
    x"05",
    x"32",
    x"28",
    x"e0",
    x"3a",
    x"63",
    x"e0",
    x"32",
    x"60",
    x"e0",
    x"c3",
    x"4b",
    x"53",
    x"21",
    x"a7",
    x"e0",
    x"5e",
    x"4b",
    x"16",
    x"e3",
    x"eb",
    x"7e",
    x"a7",
    x"c2",
    x"6f",
    x"53",
    x"1b",
    x"1a",
    x"6f",
    x"26",
    x"e4",
    x"7e",
    x"fe",
    x"02",
    x"20",
    x"30",
    x"7d",
    x"c6",
    x"09",
    x"6f",
    x"7e",
    x"b9",
    x"20",
    x"28",
    x"af",
    x"32",
    x"a5",
    x"e0",
    x"1a",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"c6",
    x"80",
    x"6f",
    x"26",
    x"e7",
    x"11",
    x"b0",
    x"e7",
    x"7e",
    x"2c",
    x"d6",
    x"10",
    x"12",
    x"1c",
    x"7e",
    x"2c",
    x"12",
    x"1c",
    x"7e",
    x"e6",
    x"1f",
    x"12",
    x"c3",
    x"6f",
    x"53",
    x"7d",
    x"e6",
    x"f0",
    x"12",
    x"18",
    x"d8",
    x"21",
    x"00",
    x"e4",
    x"06",
    x"0c",
    x"7e",
    x"fe",
    x"02",
    x"28",
    x"08",
    x"7d",
    x"c6",
    x"10",
    x"6f",
    x"10",
    x"f5",
    x"18",
    x"0f",
    x"7d",
    x"c6",
    x"09",
    x"6f",
    x"7e",
    x"b9",
    x"ca",
    x"c1",
    x"56",
    x"7d",
    x"c6",
    x"07",
    x"6f",
    x"10",
    x"e4",
    x"21",
    x"b0",
    x"e7",
    x"7e",
    x"3c",
    x"c2",
    x"3e",
    x"55",
    x"2c",
    x"2c",
    x"7e",
    x"a7",
    x"c2",
    x"3e",
    x"55",
    x"3e",
    x"06",
    x"32",
    x"28",
    x"e0",
    x"3e",
    x"01",
    x"32",
    x"a5",
    x"e0",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"c3",
    x"6f",
    x"53",
    x"cd",
    x"6e",
    x"41",
    x"3a",
    x"b4",
    x"e7",
    x"d6",
    x"80",
    x"fe",
    x"28",
    x"d2",
    x"d3",
    x"57",
    x"3a",
    x"28",
    x"e0",
    x"fe",
    x"03",
    x"ca",
    x"d3",
    x"57",
    x"21",
    x"21",
    x"e0",
    x"7e",
    x"a7",
    x"20",
    x"10",
    x"23",
    x"7e",
    x"a7",
    x"ca",
    x"d3",
    x"57",
    x"21",
    x"25",
    x"e0",
    x"34",
    x"7e",
    x"fe",
    x"14",
    x"da",
    x"d3",
    x"57",
    x"af",
    x"32",
    x"25",
    x"e0",
    x"21",
    x"30",
    x"e1",
    x"11",
    x"06",
    x"00",
    x"06",
    x"02",
    x"cb",
    x"7e",
    x"28",
    x"06",
    x"19",
    x"10",
    x"f9",
    x"c3",
    x"d3",
    x"57",
    x"3e",
    x"01",
    x"32",
    x"90",
    x"e1",
    x"ed",
    x"5b",
    x"f0",
    x"e0",
    x"13",
    x"ed",
    x"53",
    x"f0",
    x"e0",
    x"3a",
    x"28",
    x"e0",
    x"3d",
    x"ca",
    x"aa",
    x"57",
    x"36",
    x"80",
    x"23",
    x"3a",
    x"b6",
    x"e7",
    x"4f",
    x"0f",
    x"11",
    x"9a",
    x"57",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"13",
    x"77",
    x"23",
    x"36",
    x"00",
    x"23",
    x"1a",
    x"77",
    x"23",
    x"36",
    x"00",
    x"21",
    x"b8",
    x"e7",
    x"05",
    x"20",
    x"04",
    x"7d",
    x"c6",
    x"04",
    x"6f",
    x"11",
    x"b4",
    x"e7",
    x"1a",
    x"1c",
    x"77",
    x"2c",
    x"1a",
    x"1c",
    x"77",
    x"2c",
    x"1a",
    x"c6",
    x"b0",
    x"77",
    x"2c",
    x"36",
    x"0f",
    x"c3",
    x"d3",
    x"57",
    x"b3",
    x"00",
    x"bf",
    x"41",
    x"00",
    x"4d",
    x"41",
    x"41",
    x"4d",
    x"00",
    x"41",
    x"bf",
    x"00",
    x"b3",
    x"bf",
    x"bf",
    x"36",
    x"81",
    x"23",
    x"36",
    x"b3",
    x"23",
    x"af",
    x"77",
    x"23",
    x"77",
    x"23",
    x"77",
    x"21",
    x"b8",
    x"e7",
    x"05",
    x"20",
    x"04",
    x"7d",
    x"c6",
    x"04",
    x"6f",
    x"11",
    x"b4",
    x"e7",
    x"1a",
    x"1c",
    x"77",
    x"2c",
    x"1a",
    x"1c",
    x"c6",
    x"06",
    x"77",
    x"2c",
    x"3e",
    x"d0",
    x"77",
    x"2c",
    x"36",
    x"0f",
    x"21",
    x"30",
    x"e1",
    x"11",
    x"b8",
    x"e7",
    x"06",
    x"02",
    x"e5",
    x"d5",
    x"cb",
    x"7e",
    x"ca",
    x"14",
    x"58",
    x"23",
    x"7e",
    x"23",
    x"cd",
    x"26",
    x"58",
    x"4f",
    x"1a",
    x"81",
    x"12",
    x"fe",
    x"f8",
    x"30",
    x"04",
    x"fe",
    x"b8",
    x"30",
    x"10",
    x"13",
    x"23",
    x"7e",
    x"23",
    x"cd",
    x"26",
    x"58",
    x"4f",
    x"1a",
    x"81",
    x"12",
    x"fe",
    x"ba",
    x"da",
    x"14",
    x"58",
    x"2a",
    x"f2",
    x"e0",
    x"23",
    x"22",
    x"f2",
    x"e0",
    x"3e",
    x"e0",
    x"d1",
    x"12",
    x"e1",
    x"36",
    x"00",
    x"18",
    x"02",
    x"d1",
    x"e1",
    x"7b",
    x"c6",
    x"04",
    x"5f",
    x"3e",
    x"06",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"10",
    x"b8",
    x"c3",
    x"08",
    x"57",
    x"86",
    x"fa",
    x"36",
    x"58",
    x"4f",
    x"e6",
    x"0f",
    x"77",
    x"79",
    x"e6",
    x"f0",
    x"1f",
    x"1f",
    x"1f",
    x"1f",
    x"c9",
    x"4f",
    x"f6",
    x"f0",
    x"77",
    x"79",
    x"2f",
    x"e6",
    x"f0",
    x"1f",
    x"1f",
    x"1f",
    x"1f",
    x"ed",
    x"44",
    x"c9",
    x"cd",
    x"6e",
    x"41",
    x"3a",
    x"0d",
    x"e0",
    x"3d",
    x"28",
    x"08",
    x"3a",
    x"09",
    x"e0",
    x"e6",
    x"01",
    x"ca",
    x"fa",
    x"58",
    x"21",
    x"1a",
    x"e0",
    x"7e",
    x"a7",
    x"28",
    x"04",
    x"35",
    x"c3",
    x"fa",
    x"58",
    x"3a",
    x"18",
    x"e0",
    x"a7",
    x"c2",
    x"fa",
    x"58",
    x"3a",
    x"80",
    x"e0",
    x"47",
    x"21",
    x"92",
    x"e0",
    x"7e",
    x"b8",
    x"d2",
    x"fa",
    x"58",
    x"21",
    x"a4",
    x"e0",
    x"7e",
    x"fe",
    x"30",
    x"38",
    x"02",
    x"3e",
    x"fc",
    x"c6",
    x"04",
    x"77",
    x"47",
    x"11",
    x"80",
    x"e7",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"3a",
    x"70",
    x"e0",
    x"e6",
    x"3c",
    x"0f",
    x"0f",
    x"c6",
    x"50",
    x"67",
    x"1a",
    x"bc",
    x"d2",
    x"fa",
    x"58",
    x"21",
    x"04",
    x"e4",
    x"78",
    x"87",
    x"87",
    x"85",
    x"6f",
    x"7e",
    x"e6",
    x"7f",
    x"c2",
    x"fa",
    x"58",
    x"2c",
    x"7e",
    x"97",
    x"fe",
    x"0b",
    x"30",
    x"4c",
    x"7d",
    x"c6",
    x"06",
    x"6f",
    x"7e",
    x"3d",
    x"fa",
    x"fa",
    x"58",
    x"77",
    x"21",
    x"92",
    x"e0",
    x"34",
    x"21",
    x"40",
    x"e1",
    x"7e",
    x"a7",
    x"28",
    x"06",
    x"2c",
    x"2c",
    x"2c",
    x"2c",
    x"18",
    x"f6",
    x"36",
    x"01",
    x"e5",
    x"01",
    x"80",
    x"06",
    x"09",
    x"1a",
    x"47",
    x"1c",
    x"77",
    x"2c",
    x"1a",
    x"4f",
    x"77",
    x"2c",
    x"e5",
    x"50",
    x"59",
    x"cd",
    x"8a",
    x"59",
    x"fe",
    x"12",
    x"20",
    x"02",
    x"3e",
    x"11",
    x"fe",
    x"00",
    x"20",
    x"02",
    x"3e",
    x"0e",
    x"4f",
    x"e1",
    x"36",
    x"c0",
    x"2c",
    x"36",
    x"0e",
    x"e1",
    x"2c",
    x"71",
    x"2c",
    x"af",
    x"77",
    x"2c",
    x"77",
    x"21",
    x"40",
    x"e1",
    x"dd",
    x"21",
    x"c0",
    x"e7",
    x"06",
    x"08",
    x"c5",
    x"7e",
    x"a7",
    x"28",
    x"05",
    x"e5",
    x"cd",
    x"19",
    x"59",
    x"e1",
    x"01",
    x"04",
    x"00",
    x"09",
    x"dd",
    x"09",
    x"c1",
    x"10",
    x"ed",
    x"c3",
    x"45",
    x"58",
    x"23",
    x"7e",
    x"4f",
    x"23",
    x"11",
    x"c0",
    x"9f",
    x"83",
    x"5f",
    x"1a",
    x"86",
    x"c6",
    x"08",
    x"47",
    x"fa",
    x"32",
    x"59",
    x"fe",
    x"10",
    x"38",
    x"15",
    x"e6",
    x"f0",
    x"18",
    x"02",
    x"f6",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"dd",
    x"86",
    x"00",
    x"fe",
    x"c0",
    x"d2",
    x"7d",
    x"59",
    x"dd",
    x"77",
    x"00",
    x"78",
    x"e6",
    x"0f",
    x"d6",
    x"08",
    x"77",
    x"23",
    x"7b",
    x"c6",
    x"08",
    x"e6",
    x"1f",
    x"47",
    x"7b",
    x"e6",
    x"e0",
    x"b0",
    x"5f",
    x"1a",
    x"86",
    x"c6",
    x"08",
    x"47",
    x"fa",
    x"65",
    x"59",
    x"fe",
    x"10",
    x"38",
    x"14",
    x"e6",
    x"f0",
    x"18",
    x"02",
    x"f6",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"dd",
    x"86",
    x"01",
    x"dd",
    x"77",
    x"01",
    x"fe",
    x"bc",
    x"30",
    x"07",
    x"78",
    x"e6",
    x"0f",
    x"d6",
    x"08",
    x"77",
    x"c9",
    x"2d",
    x"2d",
    x"2d",
    x"36",
    x"00",
    x"dd",
    x"36",
    x"00",
    x"e0",
    x"21",
    x"92",
    x"e0",
    x"35",
    x"c9",
    x"c5",
    x"21",
    x"b4",
    x"e7",
    x"7e",
    x"2c",
    x"6e",
    x"67",
    x"3a",
    x"28",
    x"e0",
    x"3d",
    x"20",
    x"04",
    x"7d",
    x"c6",
    x"07",
    x"6f",
    x"eb",
    x"cd",
    x"d4",
    x"52",
    x"c1",
    x"fe",
    x"0d",
    x"30",
    x"02",
    x"3e",
    x"0d",
    x"fe",
    x"13",
    x"d8",
    x"3e",
    x"12",
    x"c9",
    x"cd",
    x"a1",
    x"8a",
    x"cd",
    x"e5",
    x"89",
    x"cd",
    x"9c",
    x"95",
    x"cd",
    x"ae",
    x"98",
    x"cd",
    x"7d",
    x"41",
    x"cd",
    x"c4",
    x"59",
    x"21",
    x"02",
    x"e0",
    x"36",
    x"03",
    x"06",
    x"1e",
    x"cd",
    x"c2",
    x"8a",
    x"10",
    x"fb",
    x"21",
    x"01",
    x"ef",
    x"06",
    x"18",
    x"cd",
    x"c2",
    x"8a",
    x"e6",
    x"03",
    x"c6",
    x"20",
    x"cb",
    x"40",
    x"28",
    x"02",
    x"c6",
    x"04",
    x"77",
    x"2c",
    x"10",
    x"ef",
    x"21",
    x"01",
    x"ef",
    x"11",
    x"21",
    x"ef",
    x"06",
    x"df",
    x"c5",
    x"7e",
    x"a7",
    x"28",
    x"09",
    x"47",
    x"e6",
    x"fc",
    x"4f",
    x"04",
    x"78",
    x"e6",
    x"03",
    x"b1",
    x"12",
    x"1c",
    x"2c",
    x"c1",
    x"10",
    x"ec",
    x"06",
    x"18",
    x"cd",
    x"c2",
    x"8a",
    x"6f",
    x"e6",
    x"03",
    x"c6",
    x"03",
    x"4f",
    x"7d",
    x"e6",
    x"e0",
    x"80",
    x"6f",
    x"36",
    x"00",
    x"c6",
    x"20",
    x"6f",
    x"0d",
    x"20",
    x"f8",
    x"10",
    x"e8",
    x"21",
    x"01",
    x"ef",
    x"70",
    x"2c",
    x"70",
    x"c9",
    x"21",
    x"00",
    x"e1",
    x"06",
    x"01",
    x"cd",
    x"e1",
    x"8a",
    x"af",
    x"32",
    x"28",
    x"e0",
    x"32",
    x"a8",
    x"e0",
    x"af",
    x"32",
    x"45",
    x"e0",
    x"3e",
    x"03",
    x"32",
    x"47",
    x"e0",
    x"3e",
    x"07",
    x"32",
    x"48",
    x"e0",
    x"3e",
    x"ff",
    x"32",
    x"46",
    x"e0",
    x"21",
    x"40",
    x"e0",
    x"af",
    x"06",
    x"04",
    x"77",
    x"23",
    x"10",
    x"fc",
    x"3e",
    x"01",
    x"32",
    x"44",
    x"e0",
    x"01",
    x"00",
    x"00",
    x"ed",
    x"43",
    x"70",
    x"e0",
    x"ed",
    x"43",
    x"72",
    x"e0",
    x"af",
    x"32",
    x"75",
    x"e0",
    x"3e",
    x"03",
    x"32",
    x"0e",
    x"e0",
    x"cd",
    x"79",
    x"5a",
    x"cd",
    x"e8",
    x"5a",
    x"21",
    x"75",
    x"5a",
    x"11",
    x"58",
    x"e0",
    x"01",
    x"04",
    x"00",
    x"ed",
    x"b0",
    x"c9",
    x"06",
    x"0c",
    x"09",
    x"05",
    x"af",
    x"21",
    x"14",
    x"e0",
    x"77",
    x"23",
    x"77",
    x"23",
    x"77",
    x"21",
    x"30",
    x"e3",
    x"06",
    x"03",
    x"cd",
    x"e1",
    x"8a",
    x"11",
    x"2d",
    x"e3",
    x"21",
    x"dc",
    x"5a",
    x"01",
    x"04",
    x"00",
    x"ed",
    x"b0",
    x"21",
    x"32",
    x"e3",
    x"0e",
    x"04",
    x"3e",
    x"1d",
    x"06",
    x"0a",
    x"77",
    x"23",
    x"c6",
    x"0f",
    x"10",
    x"fa",
    x"0d",
    x"20",
    x"f3",
    x"3e",
    x"0f",
    x"06",
    x"04",
    x"21",
    x"5a",
    x"e3",
    x"77",
    x"23",
    x"10",
    x"fc",
    x"36",
    x"ff",
    x"21",
    x"51",
    x"e0",
    x"36",
    x"ff",
    x"23",
    x"36",
    x"00",
    x"21",
    x"10",
    x"e0",
    x"36",
    x"28",
    x"23",
    x"36",
    x"04",
    x"23",
    x"36",
    x"10",
    x"23",
    x"36",
    x"14",
    x"11",
    x"89",
    x"e3",
    x"21",
    x"e0",
    x"5a",
    x"0e",
    x"08",
    x"ed",
    x"b0",
    x"21",
    x"c0",
    x"e8",
    x"06",
    x"0c",
    x"c3",
    x"e1",
    x"8a",
    x"48",
    x"58",
    x"68",
    x"78",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"00",
    x"03",
    x"00",
    x"21",
    x"b0",
    x"e7",
    x"36",
    x"e0",
    x"23",
    x"36",
    x"75",
    x"23",
    x"36",
    x"00",
    x"23",
    x"36",
    x"0f",
    x"c9",
    x"af",
    x"32",
    x"d4",
    x"e4",
    x"32",
    x"dc",
    x"e4",
    x"32",
    x"d7",
    x"e4",
    x"32",
    x"91",
    x"e0",
    x"32",
    x"a0",
    x"e0",
    x"32",
    x"a1",
    x"e0",
    x"21",
    x"8c",
    x"e0",
    x"77",
    x"23",
    x"77",
    x"3c",
    x"32",
    x"0d",
    x"e0",
    x"21",
    x"8e",
    x"e0",
    x"77",
    x"2c",
    x"36",
    x"18",
    x"2c",
    x"36",
    x"20",
    x"21",
    x"75",
    x"e0",
    x"7e",
    x"4f",
    x"3c",
    x"fe",
    x"1b",
    x"38",
    x"02",
    x"3e",
    x"17",
    x"77",
    x"79",
    x"3c",
    x"3c",
    x"e6",
    x"03",
    x"ca",
    x"85",
    x"5c",
    x"79",
    x"3c",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"ed",
    x"44",
    x"81",
    x"87",
    x"4f",
    x"87",
    x"81",
    x"21",
    x"0d",
    x"5c",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"79",
    x"32",
    x"8b",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"4f",
    x"e6",
    x"0e",
    x"0f",
    x"eb",
    x"21",
    x"07",
    x"5c",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"22",
    x"d0",
    x"e4",
    x"eb",
    x"79",
    x"e6",
    x"01",
    x"32",
    x"dd",
    x"e4",
    x"78",
    x"32",
    x"d5",
    x"e4",
    x"cd",
    x"f7",
    x"5b",
    x"4f",
    x"87",
    x"81",
    x"32",
    x"87",
    x"e0",
    x"78",
    x"87",
    x"80",
    x"32",
    x"89",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"87",
    x"87",
    x"32",
    x"94",
    x"e0",
    x"78",
    x"87",
    x"80",
    x"32",
    x"83",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"4f",
    x"e6",
    x"08",
    x"32",
    x"85",
    x"e0",
    x"79",
    x"e6",
    x"07",
    x"32",
    x"23",
    x"e1",
    x"78",
    x"32",
    x"84",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"32",
    x"95",
    x"e0",
    x"78",
    x"32",
    x"96",
    x"e0",
    x"cd",
    x"f7",
    x"5b",
    x"32",
    x"aa",
    x"e0",
    x"78",
    x"32",
    x"60",
    x"e0",
    x"32",
    x"63",
    x"e0",
    x"3a",
    x"75",
    x"e0",
    x"3c",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"3d",
    x"fe",
    x"03",
    x"38",
    x"04",
    x"d6",
    x"03",
    x"18",
    x"f8",
    x"47",
    x"87",
    x"80",
    x"87",
    x"21",
    x"e5",
    x"5b",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"78",
    x"11",
    x"98",
    x"e0",
    x"01",
    x"06",
    x"00",
    x"ed",
    x"b0",
    x"cd",
    x"c6",
    x"95",
    x"21",
    x"b8",
    x"4c",
    x"22",
    x"9e",
    x"e0",
    x"c9",
    x"6d",
    x"8c",
    x"93",
    x"8c",
    x"96",
    x"8c",
    x"ab",
    x"8c",
    x"cf",
    x"8c",
    x"e2",
    x"8c",
    x"f2",
    x"8c",
    x"15",
    x"8d",
    x"2b",
    x"8d",
    x"7e",
    x"23",
    x"47",
    x"e6",
    x"f0",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"08",
    x"78",
    x"e6",
    x"0f",
    x"47",
    x"08",
    x"c9",
    x"36",
    x"4c",
    x"5e",
    x"4c",
    x"86",
    x"4c",
    x"40",
    x"00",
    x"00",
    x"46",
    x"00",
    x"04",
    x"80",
    x"11",
    x"00",
    x"47",
    x"20",
    x"04",
    x"01",
    x"21",
    x"11",
    x"37",
    x"21",
    x"b5",
    x"81",
    x"32",
    x"11",
    x"38",
    x"21",
    x"b5",
    x"41",
    x"42",
    x"21",
    x"38",
    x"21",
    x"b5",
    x"11",
    x"52",
    x"22",
    x"b9",
    x"21",
    x"d6",
    x"92",
    x"63",
    x"22",
    x"a9",
    x"31",
    x"d6",
    x"40",
    x"11",
    x"10",
    x"b7",
    x"01",
    x"d6",
    x"12",
    x"64",
    x"32",
    x"a7",
    x"31",
    x"e7",
    x"93",
    x"76",
    x"32",
    x"a8",
    x"41",
    x"e7",
    x"53",
    x"76",
    x"32",
    x"a8",
    x"41",
    x"e7",
    x"13",
    x"87",
    x"42",
    x"a9",
    x"41",
    x"b8",
    x"94",
    x"87",
    x"42",
    x"a9",
    x"61",
    x"b8",
    x"50",
    x"22",
    x"11",
    x"b7",
    x"21",
    x"b8",
    x"13",
    x"88",
    x"52",
    x"9a",
    x"61",
    x"d8",
    x"94",
    x"88",
    x"52",
    x"9a",
    x"61",
    x"d8",
    x"54",
    x"88",
    x"52",
    x"9c",
    x"61",
    x"d8",
    x"13",
    x"98",
    x"62",
    x"9c",
    x"71",
    x"e8",
    x"94",
    x"99",
    x"62",
    x"9c",
    x"71",
    x"e8",
    x"54",
    x"99",
    x"62",
    x"9c",
    x"71",
    x"e8",
    x"21",
    x"0d",
    x"e0",
    x"36",
    x"03",
    x"3e",
    x"1e",
    x"32",
    x"a2",
    x"e0",
    x"3a",
    x"71",
    x"e0",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"4f",
    x"e6",
    x"07",
    x"47",
    x"21",
    x"cf",
    x"5c",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"c5",
    x"cd",
    x"c6",
    x"95",
    x"c1",
    x"78",
    x"87",
    x"21",
    x"0b",
    x"5d",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"22",
    x"d0",
    x"e4",
    x"21",
    x"d7",
    x"5c",
    x"22",
    x"9e",
    x"e0",
    x"79",
    x"fe",
    x"06",
    x"3e",
    x"03",
    x"30",
    x"03",
    x"78",
    x"cb",
    x"3f",
    x"c6",
    x"0b",
    x"32",
    x"aa",
    x"e0",
    x"c9",
    x"05",
    x"06",
    x"03",
    x"00",
    x"07",
    x"01",
    x"02",
    x"04",
    x"ff",
    x"fc",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"ff",
    x"f1",
    x"c0",
    x"00",
    x"c0",
    x"00",
    x"c0",
    x"00",
    x"c0",
    x"00",
    x"ff",
    x"f1",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"ff",
    x"f0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"ff",
    x"f0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"ff",
    x"fe",
    x"1b",
    x"5d",
    x"43",
    x"5d",
    x"6b",
    x"5d",
    x"93",
    x"5d",
    x"bb",
    x"5d",
    x"e3",
    x"5d",
    x"0b",
    x"5e",
    x"33",
    x"5e",
    x"08",
    x"00",
    x"40",
    x"8d",
    x"00",
    x"40",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"52",
    x"8d",
    x"00",
    x"52",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"52",
    x"8d",
    x"80",
    x"52",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"40",
    x"8d",
    x"00",
    x"40",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"40",
    x"8d",
    x"80",
    x"40",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"6a",
    x"8d",
    x"00",
    x"6a",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"81",
    x"8d",
    x"00",
    x"81",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"81",
    x"8d",
    x"00",
    x"81",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"6a",
    x"8d",
    x"00",
    x"6a",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"6a",
    x"8d",
    x"80",
    x"6a",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"91",
    x"8d",
    x"00",
    x"a8",
    x"8d",
    x"00",
    x"08",
    x"00",
    x"bf",
    x"8d",
    x"00",
    x"bf",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"bf",
    x"8d",
    x"00",
    x"bf",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"91",
    x"8d",
    x"00",
    x"a8",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"91",
    x"8d",
    x"80",
    x"a8",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"e0",
    x"8d",
    x"00",
    x"db",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"fe",
    x"8d",
    x"00",
    x"fe",
    x"8d",
    x"00",
    x"08",
    x"08",
    x"fe",
    x"8d",
    x"80",
    x"fe",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"e0",
    x"8d",
    x"00",
    x"db",
    x"8d",
    x"80",
    x"08",
    x"00",
    x"db",
    x"8d",
    x"00",
    x"e0",
    x"8d",
    x"80",
    x"08",
    x"08",
    x"2f",
    x"8e",
    x"00",
    x"2f",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"57",
    x"8e",
    x"00",
    x"57",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"57",
    x"8e",
    x"80",
    x"57",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"2f",
    x"8e",
    x"00",
    x"2f",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"2f",
    x"8e",
    x"80",
    x"2f",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"7a",
    x"8e",
    x"00",
    x"7a",
    x"8e",
    x"00",
    x"08",
    x"00",
    x"9f",
    x"8e",
    x"00",
    x"9f",
    x"8e",
    x"80",
    x"08",
    x"00",
    x"9f",
    x"8e",
    x"00",
    x"9f",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"7a",
    x"8e",
    x"00",
    x"7a",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"7a",
    x"8e",
    x"80",
    x"7a",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"bd",
    x"8e",
    x"00",
    x"bd",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"d9",
    x"8e",
    x"00",
    x"d9",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"d9",
    x"8e",
    x"80",
    x"d9",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"bd",
    x"8e",
    x"00",
    x"bd",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"bd",
    x"8e",
    x"80",
    x"bd",
    x"8e",
    x"80",
    x"08",
    x"08",
    x"f5",
    x"8e",
    x"00",
    x"f5",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"09",
    x"8f",
    x"00",
    x"09",
    x"8f",
    x"00",
    x"08",
    x"08",
    x"09",
    x"8f",
    x"80",
    x"09",
    x"8f",
    x"80",
    x"08",
    x"08",
    x"f5",
    x"8e",
    x"00",
    x"f5",
    x"8e",
    x"00",
    x"08",
    x"08",
    x"f5",
    x"8e",
    x"80",
    x"f5",
    x"8e",
    x"80",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"8c",
    x"e0",
    x"7e",
    x"3c",
    x"fe",
    x"3c",
    x"38",
    x"09",
    x"23",
    x"7e",
    x"3c",
    x"20",
    x"01",
    x"3d",
    x"77",
    x"af",
    x"2b",
    x"77",
    x"23",
    x"4e",
    x"79",
    x"06",
    x"00",
    x"fe",
    x"1e",
    x"38",
    x"06",
    x"04",
    x"fe",
    x"3c",
    x"38",
    x"01",
    x"04",
    x"11",
    x"87",
    x"e0",
    x"21",
    x"0f",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"11",
    x"89",
    x"e0",
    x"21",
    x"2d",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"79",
    x"06",
    x"00",
    x"fe",
    x"28",
    x"38",
    x"01",
    x"04",
    x"11",
    x"8b",
    x"e0",
    x"21",
    x"4b",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"3a",
    x"10",
    x"e0",
    x"06",
    x"00",
    x"fe",
    x"14",
    x"30",
    x"09",
    x"04",
    x"04",
    x"fe",
    x"0a",
    x"30",
    x"08",
    x"04",
    x"18",
    x"05",
    x"fe",
    x"1e",
    x"30",
    x"01",
    x"04",
    x"11",
    x"94",
    x"e0",
    x"21",
    x"73",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"3a",
    x"0d",
    x"e0",
    x"3d",
    x"3e",
    x"08",
    x"20",
    x"03",
    x"3a",
    x"95",
    x"e0",
    x"32",
    x"80",
    x"e0",
    x"05",
    x"f2",
    x"d7",
    x"5e",
    x"06",
    x"00",
    x"11",
    x"83",
    x"e0",
    x"21",
    x"93",
    x"5f",
    x"cd",
    x"04",
    x"5f",
    x"3a",
    x"17",
    x"e0",
    x"a7",
    x"c2",
    x"5b",
    x"5e",
    x"21",
    x"10",
    x"e0",
    x"3a",
    x"84",
    x"e0",
    x"be",
    x"da",
    x"5b",
    x"5e",
    x"21",
    x"0d",
    x"e0",
    x"7e",
    x"3d",
    x"ca",
    x"5b",
    x"5e",
    x"3e",
    x"02",
    x"77",
    x"3e",
    x"07",
    x"32",
    x"8a",
    x"e0",
    x"c3",
    x"5b",
    x"5e",
    x"1a",
    x"80",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"1b",
    x"12",
    x"c9",
    x"60",
    x"50",
    x"40",
    x"50",
    x"40",
    x"30",
    x"50",
    x"30",
    x"30",
    x"40",
    x"30",
    x"20",
    x"40",
    x"20",
    x"20",
    x"30",
    x"30",
    x"20",
    x"30",
    x"20",
    x"10",
    x"20",
    x"20",
    x"10",
    x"20",
    x"10",
    x"10",
    x"10",
    x"10",
    x"10",
    x"90",
    x"70",
    x"50",
    x"80",
    x"60",
    x"40",
    x"70",
    x"50",
    x"40",
    x"60",
    x"40",
    x"30",
    x"50",
    x"30",
    x"30",
    x"40",
    x"30",
    x"30",
    x"40",
    x"20",
    x"20",
    x"30",
    x"30",
    x"20",
    x"30",
    x"20",
    x"20",
    x"20",
    x"20",
    x"20",
    x"02",
    x"02",
    x"02",
    x"03",
    x"02",
    x"03",
    x"02",
    x"03",
    x"03",
    x"03",
    x"03",
    x"03",
    x"03",
    x"04",
    x"02",
    x"03",
    x"03",
    x"04",
    x"04",
    x"04",
    x"04",
    x"05",
    x"04",
    x"05",
    x"04",
    x"05",
    x"02",
    x"03",
    x"04",
    x"06",
    x"05",
    x"06",
    x"05",
    x"06",
    x"05",
    x"07",
    x"05",
    x"07",
    x"05",
    x"07",
    x"01",
    x"01",
    x"02",
    x"02",
    x"01",
    x"02",
    x"02",
    x"02",
    x"01",
    x"02",
    x"02",
    x"03",
    x"02",
    x"02",
    x"02",
    x"03",
    x"02",
    x"02",
    x"03",
    x"03",
    x"02",
    x"02",
    x"03",
    x"04",
    x"02",
    x"03",
    x"03",
    x"04",
    x"03",
    x"03",
    x"03",
    x"04",
    x"07",
    x"05",
    x"03",
    x"06",
    x"04",
    x"02",
    x"05",
    x"03",
    x"02",
    x"89",
    x"08",
    x"86",
    x"08",
    x"87",
    x"70",
    x"88",
    x"02",
    x"03",
    x"03",
    x"c7",
    x"48",
    x"c9",
    x"04",
    x"8a",
    x"c8",
    x"04",
    x"82",
    x"ee",
    x"5f",
    x"89",
    x"08",
    x"86",
    x"08",
    x"87",
    x"80",
    x"88",
    x"02",
    x"03",
    x"03",
    x"58",
    x"58",
    x"80",
    x"58",
    x"c9",
    x"07",
    x"81",
    x"8a",
    x"c8",
    x"07",
    x"82",
    x"ee",
    x"5f",
    x"89",
    x"0f",
    x"86",
    x"50",
    x"87",
    x"f1",
    x"88",
    x"02",
    x"50",
    x"c2",
    x"06",
    x"0a",
    x"c4",
    x"50",
    x"8a",
    x"cb",
    x"27",
    x"82",
    x"ee",
    x"5f",
    x"89",
    x"0f",
    x"86",
    x"40",
    x"87",
    x"f1",
    x"88",
    x"02",
    x"58",
    x"c3",
    x"06",
    x"c5",
    x"4f",
    x"8a",
    x"cc",
    x"24",
    x"82",
    x"ee",
    x"5f",
    x"84",
    x"02",
    x"85",
    x"00",
    x"84",
    x"01",
    x"84",
    x"03",
    x"84",
    x"05",
    x"84",
    x"0e",
    x"1e",
    x"88",
    x"01",
    x"82",
    x"ee",
    x"5f",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"74",
    x"e0",
    x"7e",
    x"a7",
    x"28",
    x"f6",
    x"fe",
    x"ff",
    x"28",
    x"0c",
    x"3d",
    x"77",
    x"20",
    x"ee",
    x"21",
    x"75",
    x"81",
    x"cd",
    x"8f",
    x"8a",
    x"18",
    x"e6",
    x"36",
    x"78",
    x"06",
    x"3c",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"c1",
    x"10",
    x"f9",
    x"cd",
    x"de",
    x"80",
    x"21",
    x"71",
    x"e0",
    x"34",
    x"20",
    x"03",
    x"2b",
    x"34",
    x"23",
    x"4e",
    x"23",
    x"23",
    x"7e",
    x"c6",
    x"01",
    x"27",
    x"77",
    x"2b",
    x"7e",
    x"ce",
    x"00",
    x"27",
    x"77",
    x"79",
    x"3c",
    x"e6",
    x"03",
    x"28",
    x"14",
    x"21",
    x"6d",
    x"81",
    x"cd",
    x"7e",
    x"8a",
    x"21",
    x"8e",
    x"19",
    x"11",
    x"72",
    x"e0",
    x"01",
    x"03",
    x"02",
    x"cd",
    x"4f",
    x"8a",
    x"18",
    x"16",
    x"3e",
    x"01",
    x"32",
    x"68",
    x"e2",
    x"32",
    x"70",
    x"e2",
    x"32",
    x"78",
    x"e2",
    x"21",
    x"75",
    x"81",
    x"cd",
    x"7e",
    x"8a",
    x"3e",
    x"78",
    x"32",
    x"74",
    x"e0",
    x"3a",
    x"71",
    x"e0",
    x"4f",
    x"21",
    x"19",
    x"1a",
    x"06",
    x"06",
    x"11",
    x"55",
    x"81",
    x"78",
    x"3d",
    x"87",
    x"87",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"b9",
    x"38",
    x"07",
    x"28",
    x"05",
    x"10",
    x"ec",
    x"c3",
    x"00",
    x"80",
    x"91",
    x"ed",
    x"44",
    x"4f",
    x"3e",
    x"01",
    x"32",
    x"80",
    x"e2",
    x"13",
    x"1a",
    x"47",
    x"85",
    x"e6",
    x"10",
    x"20",
    x"08",
    x"7d",
    x"e6",
    x"e0",
    x"f6",
    x"19",
    x"c6",
    x"40",
    x"6f",
    x"e5",
    x"cd",
    x"be",
    x"80",
    x"e1",
    x"7d",
    x"80",
    x"6f",
    x"06",
    x"08",
    x"e5",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"c1",
    x"10",
    x"f9",
    x"e1",
    x"c3",
    x"76",
    x"80",
    x"cd",
    x"c1",
    x"80",
    x"13",
    x"1a",
    x"c5",
    x"e5",
    x"cd",
    x"cf",
    x"80",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"c1",
    x"c9",
    x"4f",
    x"cd",
    x"4d",
    x"00",
    x"23",
    x"0c",
    x"79",
    x"10",
    x"f8",
    x"c9",
    x"21",
    x"19",
    x"19",
    x"18",
    x"03",
    x"21",
    x"19",
    x"1a",
    x"06",
    x"08",
    x"c5",
    x"01",
    x"06",
    x"00",
    x"af",
    x"cd",
    x"56",
    x"00",
    x"7d",
    x"c6",
    x"20",
    x"6f",
    x"c1",
    x"10",
    x"f1",
    x"c9",
    x"21",
    x"0e",
    x"e0",
    x"34",
    x"20",
    x"01",
    x"35",
    x"cd",
    x"d9",
    x"80",
    x"11",
    x"0e",
    x"e0",
    x"1a",
    x"a7",
    x"c8",
    x"fe",
    x"07",
    x"30",
    x"2b",
    x"21",
    x"39",
    x"19",
    x"47",
    x"c5",
    x"e5",
    x"3e",
    x"90",
    x"06",
    x"02",
    x"cd",
    x"cf",
    x"80",
    x"e1",
    x"e5",
    x"11",
    x"20",
    x"00",
    x"19",
    x"3e",
    x"92",
    x"06",
    x"02",
    x"cd",
    x"cf",
    x"80",
    x"e1",
    x"23",
    x"23",
    x"7d",
    x"f6",
    x"e0",
    x"3c",
    x"20",
    x"04",
    x"11",
    x"5a",
    x"00",
    x"19",
    x"c1",
    x"10",
    x"da",
    x"c9",
    x"21",
    x"7c",
    x"19",
    x"01",
    x"01",
    x"01",
    x"cd",
    x"58",
    x"45",
    x"21",
    x"89",
    x"81",
    x"c3",
    x"7e",
    x"8a",
    x"21",
    x"b4",
    x"e7",
    x"36",
    x"a3",
    x"23",
    x"36",
    x"60",
    x"23",
    x"36",
    x"00",
    x"23",
    x"36",
    x"0f",
    x"21",
    x"0e",
    x"e0",
    x"35",
    x"18",
    x"a5",
    x"01",
    x"01",
    x"b4",
    x"b5",
    x"05",
    x"01",
    x"b6",
    x"b7",
    x"0a",
    x"02",
    x"b8",
    x"ba",
    x"14",
    x"02",
    x"bc",
    x"be",
    x"1e",
    x"02",
    x"c0",
    x"c2",
    x"32",
    x"02",
    x"c4",
    x"c6",
    x"89",
    x"19",
    x"05",
    x"83",
    x"84",
    x"71",
    x"77",
    x"75",
    x"85",
    x"19",
    x"11",
    x"73",
    x"78",
    x"71",
    x"7c",
    x"7c",
    x"75",
    x"7e",
    x"77",
    x"79",
    x"7e",
    x"77",
    x"00",
    x"83",
    x"84",
    x"71",
    x"77",
    x"75",
    x"5a",
    x"19",
    x"04",
    x"13",
    x"08",
    x"09",
    x"10",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"28",
    x"e0",
    x"1a",
    x"a7",
    x"20",
    x"24",
    x"3a",
    x"b4",
    x"e7",
    x"fe",
    x"a3",
    x"20",
    x"1d",
    x"21",
    x"20",
    x"e1",
    x"7e",
    x"fe",
    x"02",
    x"20",
    x"15",
    x"23",
    x"3a",
    x"b5",
    x"e7",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"fe",
    x"1e",
    x"30",
    x"08",
    x"3e",
    x"02",
    x"12",
    x"3e",
    x"01",
    x"32",
    x"18",
    x"e0",
    x"11",
    x"b8",
    x"e7",
    x"cd",
    x"e4",
    x"81",
    x"28",
    x"09",
    x"af",
    x"32",
    x"30",
    x"e1",
    x"3e",
    x"e0",
    x"32",
    x"b8",
    x"e7",
    x"11",
    x"bc",
    x"e7",
    x"cd",
    x"e4",
    x"81",
    x"ca",
    x"c3",
    x"84",
    x"af",
    x"32",
    x"36",
    x"e1",
    x"3e",
    x"e0",
    x"32",
    x"bc",
    x"e7",
    x"c3",
    x"c3",
    x"84",
    x"1a",
    x"fe",
    x"e0",
    x"c8",
    x"08",
    x"1c",
    x"1a",
    x"1d",
    x"d9",
    x"5f",
    x"08",
    x"57",
    x"3a",
    x"28",
    x"e0",
    x"3d",
    x"28",
    x"05",
    x"01",
    x"07",
    x"00",
    x"18",
    x"03",
    x"01",
    x"0f",
    x"02",
    x"21",
    x"80",
    x"e7",
    x"d9",
    x"01",
    x"00",
    x"0c",
    x"3a",
    x"28",
    x"e0",
    x"d6",
    x"05",
    x"fe",
    x"03",
    x"30",
    x"01",
    x"04",
    x"d9",
    x"7a",
    x"96",
    x"f2",
    x"17",
    x"82",
    x"ed",
    x"44",
    x"fe",
    x"06",
    x"d2",
    x"46",
    x"82",
    x"2c",
    x"7b",
    x"80",
    x"96",
    x"f2",
    x"25",
    x"82",
    x"ed",
    x"44",
    x"2d",
    x"b9",
    x"d2",
    x"46",
    x"82",
    x"7d",
    x"d9",
    x"0c",
    x"d6",
    x"80",
    x"87",
    x"87",
    x"c6",
    x"04",
    x"6f",
    x"26",
    x"e4",
    x"7e",
    x"e6",
    x"7f",
    x"32",
    x"32",
    x"e0",
    x"d6",
    x"03",
    x"fe",
    x"03",
    x"d9",
    x"38",
    x"03",
    x"cd",
    x"52",
    x"82",
    x"2c",
    x"2c",
    x"2c",
    x"2c",
    x"d9",
    x"05",
    x"c2",
    x"0f",
    x"82",
    x"c3",
    x"ac",
    x"83",
    x"d9",
    x"af",
    x"32",
    x"30",
    x"e0",
    x"7d",
    x"c6",
    x"05",
    x"6f",
    x"7e",
    x"32",
    x"31",
    x"e0",
    x"fe",
    x"2d",
    x"38",
    x"05",
    x"3e",
    x"01",
    x"32",
    x"30",
    x"e0",
    x"7d",
    x"d6",
    x"09",
    x"6f",
    x"d5",
    x"e5",
    x"7e",
    x"3d",
    x"ca",
    x"08",
    x"83",
    x"3d",
    x"ca",
    x"b2",
    x"82",
    x"3d",
    x"ca",
    x"39",
    x"83",
    x"3d",
    x"ca",
    x"46",
    x"83",
    x"3e",
    x"06",
    x"21",
    x"a9",
    x"e0",
    x"35",
    x"20",
    x"03",
    x"3a",
    x"aa",
    x"e0",
    x"32",
    x"33",
    x"e0",
    x"3e",
    x"01",
    x"32",
    x"e0",
    x"e1",
    x"3a",
    x"30",
    x"e0",
    x"a7",
    x"c2",
    x"63",
    x"83",
    x"21",
    x"10",
    x"e0",
    x"35",
    x"3a",
    x"31",
    x"e0",
    x"fe",
    x"19",
    x"30",
    x"07",
    x"21",
    x"12",
    x"e0",
    x"35",
    x"c3",
    x"63",
    x"83",
    x"21",
    x"13",
    x"e0",
    x"35",
    x"c3",
    x"63",
    x"83",
    x"d9",
    x"2c",
    x"2c",
    x"2c",
    x"7e",
    x"fe",
    x"04",
    x"28",
    x"0f",
    x"3e",
    x"01",
    x"32",
    x"f8",
    x"e1",
    x"36",
    x"04",
    x"2d",
    x"2d",
    x"2d",
    x"d9",
    x"e1",
    x"d1",
    x"d9",
    x"c9",
    x"3e",
    x"01",
    x"32",
    x"f0",
    x"e1",
    x"3e",
    x"78",
    x"32",
    x"1a",
    x"e0",
    x"2d",
    x"2d",
    x"2d",
    x"d9",
    x"3a",
    x"0d",
    x"e0",
    x"fe",
    x"03",
    x"20",
    x"0d",
    x"21",
    x"a9",
    x"e0",
    x"35",
    x"20",
    x"07",
    x"3e",
    x"ff",
    x"32",
    x"33",
    x"e0",
    x"18",
    x"0c",
    x"e5",
    x"e1",
    x"7d",
    x"c6",
    x"0c",
    x"6f",
    x"7e",
    x"c6",
    x"03",
    x"32",
    x"33",
    x"e0",
    x"e1",
    x"e5",
    x"3a",
    x"32",
    x"e0",
    x"fe",
    x"09",
    x"20",
    x"4e",
    x"3e",
    x"03",
    x"32",
    x"20",
    x"e1",
    x"18",
    x"47",
    x"af",
    x"32",
    x"a5",
    x"e0",
    x"3c",
    x"32",
    x"d0",
    x"e1",
    x"32",
    x"18",
    x"e2",
    x"32",
    x"20",
    x"e2",
    x"21",
    x"28",
    x"e0",
    x"7e",
    x"36",
    x"00",
    x"fe",
    x"05",
    x"20",
    x"04",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"21",
    x"b0",
    x"e7",
    x"7e",
    x"3c",
    x"20",
    x"04",
    x"2c",
    x"2c",
    x"7e",
    x"a7",
    x"3e",
    x"09",
    x"20",
    x"01",
    x"3d",
    x"32",
    x"33",
    x"e0",
    x"18",
    x"2a",
    x"3c",
    x"32",
    x"e8",
    x"e1",
    x"e1",
    x"e5",
    x"3e",
    x"06",
    x"32",
    x"33",
    x"e0",
    x"18",
    x"09",
    x"3c",
    x"32",
    x"e0",
    x"e1",
    x"3e",
    x"07",
    x"32",
    x"33",
    x"e0",
    x"3a",
    x"30",
    x"e0",
    x"a7",
    x"20",
    x"0e",
    x"7e",
    x"21",
    x"0f",
    x"e0",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"35",
    x"21",
    x"10",
    x"e0",
    x"35",
    x"21",
    x"a0",
    x"e0",
    x"34",
    x"21",
    x"33",
    x"e0",
    x"7e",
    x"fe",
    x"ff",
    x"20",
    x"09",
    x"3a",
    x"aa",
    x"e0",
    x"77",
    x"cd",
    x"98",
    x"85",
    x"3e",
    x"03",
    x"cd",
    x"98",
    x"85",
    x"e1",
    x"d1",
    x"36",
    x"00",
    x"d9",
    x"d5",
    x"11",
    x"d7",
    x"e4",
    x"1a",
    x"3d",
    x"12",
    x"3a",
    x"10",
    x"e1",
    x"5f",
    x"c6",
    x"04",
    x"e6",
    x"0f",
    x"32",
    x"10",
    x"e1",
    x"7b",
    x"11",
    x"00",
    x"e1",
    x"83",
    x"5f",
    x"3e",
    x"ff",
    x"12",
    x"1c",
    x"3a",
    x"33",
    x"e0",
    x"12",
    x"1c",
    x"7e",
    x"12",
    x"2c",
    x"1c",
    x"7e",
    x"12",
    x"2d",
    x"d1",
    x"36",
    x"e0",
    x"c9",
    x"d9",
    x"21",
    x"00",
    x"e3",
    x"7a",
    x"d6",
    x"0f",
    x"f2",
    x"b8",
    x"83",
    x"ed",
    x"44",
    x"fe",
    x"06",
    x"30",
    x"71",
    x"d9",
    x"06",
    x"04",
    x"d9",
    x"7e",
    x"a7",
    x"ca",
    x"28",
    x"84",
    x"e5",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7b",
    x"80",
    x"96",
    x"f2",
    x"d2",
    x"83",
    x"ed",
    x"44",
    x"b9",
    x"30",
    x"52",
    x"7d",
    x"d6",
    x"2d",
    x"6f",
    x"7e",
    x"3d",
    x"28",
    x"40",
    x"32",
    x"f0",
    x"e1",
    x"e5",
    x"21",
    x"10",
    x"e0",
    x"35",
    x"21",
    x"11",
    x"e0",
    x"35",
    x"21",
    x"14",
    x"e0",
    x"35",
    x"d5",
    x"c5",
    x"af",
    x"cd",
    x"98",
    x"85",
    x"c1",
    x"d1",
    x"e1",
    x"36",
    x"00",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"d5",
    x"3a",
    x"10",
    x"e1",
    x"5f",
    x"c6",
    x"04",
    x"e6",
    x"0f",
    x"32",
    x"10",
    x"e1",
    x"7b",
    x"11",
    x"00",
    x"e1",
    x"83",
    x"5f",
    x"3e",
    x"ff",
    x"12",
    x"1c",
    x"1c",
    x"1c",
    x"7e",
    x"12",
    x"1d",
    x"3e",
    x"0f",
    x"12",
    x"d1",
    x"18",
    x"07",
    x"36",
    x"02",
    x"3e",
    x"01",
    x"32",
    x"f8",
    x"e1",
    x"d9",
    x"0c",
    x"d9",
    x"e1",
    x"2c",
    x"d9",
    x"10",
    x"93",
    x"d9",
    x"21",
    x"5f",
    x"e3",
    x"3e",
    x"04",
    x"08",
    x"7a",
    x"96",
    x"f2",
    x"3a",
    x"84",
    x"ed",
    x"44",
    x"fe",
    x"06",
    x"d2",
    x"b6",
    x"84",
    x"e5",
    x"7d",
    x"d6",
    x"5a",
    x"6f",
    x"d9",
    x"06",
    x"0a",
    x"d9",
    x"7e",
    x"a7",
    x"28",
    x"64",
    x"e5",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7b",
    x"80",
    x"96",
    x"f2",
    x"59",
    x"84",
    x"ed",
    x"44",
    x"b9",
    x"30",
    x"53",
    x"d5",
    x"e5",
    x"08",
    x"57",
    x"08",
    x"7a",
    x"11",
    x"12",
    x"e0",
    x"21",
    x"15",
    x"e0",
    x"fe",
    x"03",
    x"30",
    x"0b",
    x"13",
    x"23",
    x"3e",
    x"01",
    x"32",
    x"e0",
    x"e1",
    x"3e",
    x"02",
    x"18",
    x"05",
    x"3e",
    x"01",
    x"32",
    x"e8",
    x"e1",
    x"35",
    x"eb",
    x"35",
    x"c5",
    x"cd",
    x"98",
    x"85",
    x"c1",
    x"21",
    x"10",
    x"e0",
    x"35",
    x"21",
    x"10",
    x"e1",
    x"7e",
    x"5e",
    x"c6",
    x"04",
    x"e6",
    x"0f",
    x"77",
    x"16",
    x"e1",
    x"e1",
    x"3e",
    x"ff",
    x"12",
    x"1c",
    x"af",
    x"12",
    x"1c",
    x"1c",
    x"7e",
    x"12",
    x"1d",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"12",
    x"d1",
    x"e1",
    x"36",
    x"00",
    x"d9",
    x"0c",
    x"d9",
    x"18",
    x"01",
    x"e1",
    x"2c",
    x"d9",
    x"10",
    x"93",
    x"d9",
    x"e1",
    x"7d",
    x"c6",
    x"0a",
    x"6f",
    x"08",
    x"3d",
    x"c2",
    x"32",
    x"84",
    x"d9",
    x"79",
    x"a7",
    x"c9",
    x"3a",
    x"28",
    x"e0",
    x"3d",
    x"fa",
    x"d9",
    x"84",
    x"28",
    x"07",
    x"fe",
    x"03",
    x"30",
    x"09",
    x"c3",
    x"90",
    x"81",
    x"21",
    x"b0",
    x"e7",
    x"cd",
    x"e2",
    x"84",
    x"21",
    x"b4",
    x"e7",
    x"cd",
    x"e2",
    x"84",
    x"c3",
    x"90",
    x"81",
    x"56",
    x"7a",
    x"fe",
    x"a3",
    x"c0",
    x"e5",
    x"2c",
    x"5e",
    x"21",
    x"80",
    x"e7",
    x"06",
    x"0c",
    x"3a",
    x"28",
    x"e0",
    x"d6",
    x"05",
    x"fe",
    x"03",
    x"30",
    x"01",
    x"04",
    x"7a",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"4f",
    x"7b",
    x"2c",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"81",
    x"38",
    x"04",
    x"fe",
    x"0e",
    x"38",
    x"26",
    x"2c",
    x"2c",
    x"2c",
    x"10",
    x"e6",
    x"21",
    x"c0",
    x"e7",
    x"06",
    x"08",
    x"7a",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"4f",
    x"7b",
    x"2c",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"81",
    x"38",
    x"04",
    x"fe",
    x"08",
    x"38",
    x"23",
    x"2c",
    x"2c",
    x"2c",
    x"10",
    x"e6",
    x"e1",
    x"c9",
    x"af",
    x"32",
    x"32",
    x"e0",
    x"2c",
    x"2c",
    x"36",
    x"04",
    x"2d",
    x"2d",
    x"2d",
    x"7d",
    x"d9",
    x"d6",
    x"80",
    x"87",
    x"87",
    x"c6",
    x"04",
    x"6f",
    x"26",
    x"e4",
    x"d9",
    x"cd",
    x"52",
    x"82",
    x"18",
    x"0d",
    x"2d",
    x"36",
    x"e0",
    x"11",
    x"80",
    x"f9",
    x"19",
    x"36",
    x"00",
    x"21",
    x"92",
    x"e0",
    x"35",
    x"e1",
    x"36",
    x"e0",
    x"11",
    x"28",
    x"e0",
    x"1a",
    x"3d",
    x"20",
    x"16",
    x"12",
    x"7d",
    x"fe",
    x"b0",
    x"ca",
    x"85",
    x"85",
    x"36",
    x"a3",
    x"2c",
    x"4e",
    x"11",
    x"b0",
    x"e7",
    x"3e",
    x"e0",
    x"12",
    x"1c",
    x"1a",
    x"77",
    x"18",
    x"0a",
    x"3e",
    x"01",
    x"32",
    x"17",
    x"e0",
    x"32",
    x"18",
    x"e0",
    x"2c",
    x"4e",
    x"21",
    x"16",
    x"e1",
    x"7e",
    x"a7",
    x"28",
    x"05",
    x"e5",
    x"cd",
    x"0a",
    x"87",
    x"e1",
    x"36",
    x"ff",
    x"23",
    x"71",
    x"c9",
    x"87",
    x"21",
    x"c7",
    x"85",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"56",
    x"23",
    x"5e",
    x"3a",
    x"0b",
    x"e0",
    x"3d",
    x"c8",
    x"3e",
    x"01",
    x"32",
    x"44",
    x"e0",
    x"21",
    x"43",
    x"e0",
    x"7e",
    x"83",
    x"27",
    x"77",
    x"2b",
    x"7e",
    x"8a",
    x"27",
    x"77",
    x"2b",
    x"7e",
    x"ce",
    x"00",
    x"27",
    x"77",
    x"2b",
    x"7e",
    x"ce",
    x"00",
    x"27",
    x"77",
    x"c9",
    x"01",
    x"50",
    x"00",
    x"80",
    x"00",
    x"50",
    x"04",
    x"00",
    x"08",
    x"00",
    x"16",
    x"00",
    x"01",
    x"60",
    x"01",
    x"00",
    x"05",
    x"00",
    x"10",
    x"00",
    x"01",
    x"60",
    x"10",
    x"00",
    x"15",
    x"00",
    x"20",
    x"00",
    x"30",
    x"00",
    x"3a",
    x"44",
    x"e0",
    x"3d",
    x"c0",
    x"32",
    x"44",
    x"e0",
    x"cd",
    x"7b",
    x"86",
    x"cd",
    x"3b",
    x"86",
    x"cd",
    x"43",
    x"86",
    x"3a",
    x"45",
    x"e0",
    x"21",
    x"46",
    x"e0",
    x"be",
    x"c8",
    x"3a",
    x"41",
    x"e0",
    x"21",
    x"47",
    x"e0",
    x"be",
    x"c0",
    x"3a",
    x"45",
    x"e0",
    x"a7",
    x"20",
    x"01",
    x"77",
    x"3c",
    x"fe",
    x"ff",
    x"28",
    x"03",
    x"32",
    x"45",
    x"e0",
    x"3a",
    x"48",
    x"e0",
    x"86",
    x"27",
    x"77",
    x"3e",
    x"01",
    x"32",
    x"a8",
    x"e1",
    x"32",
    x"b0",
    x"e1",
    x"32",
    x"10",
    x"e2",
    x"c3",
    x"f3",
    x"80",
    x"3a",
    x"09",
    x"e0",
    x"47",
    x"e6",
    x"0f",
    x"c0",
    x"21",
    x"2a",
    x"46",
    x"cb",
    x"60",
    x"c2",
    x"7e",
    x"8a",
    x"c3",
    x"8f",
    x"8a",
    x"21",
    x"59",
    x"18",
    x"11",
    x"01",
    x"e0",
    x"18",
    x"06",
    x"21",
    x"b9",
    x"18",
    x"11",
    x"40",
    x"e0",
    x"01",
    x"04",
    x"03",
    x"d5",
    x"13",
    x"cd",
    x"54",
    x"8a",
    x"d1",
    x"1a",
    x"a7",
    x"c8",
    x"fe",
    x"07",
    x"30",
    x"0e",
    x"47",
    x"11",
    x"1f",
    x"00",
    x"19",
    x"3e",
    x"3a",
    x"cd",
    x"4d",
    x"00",
    x"2b",
    x"10",
    x"f8",
    x"c9",
    x"11",
    x"1a",
    x"18",
    x"19",
    x"eb",
    x"21",
    x"75",
    x"86",
    x"01",
    x"06",
    x"00",
    x"c3",
    x"5c",
    x"00",
    x"20",
    x"47",
    x"52",
    x"45",
    x"41",
    x"54",
    x"11",
    x"40",
    x"e0",
    x"21",
    x"01",
    x"e0",
    x"06",
    x"04",
    x"1a",
    x"be",
    x"d8",
    x"20",
    x"05",
    x"1c",
    x"2c",
    x"10",
    x"f7",
    x"c9",
    x"1a",
    x"77",
    x"1c",
    x"2c",
    x"10",
    x"fa",
    x"c9",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"16",
    x"e1",
    x"7e",
    x"a7",
    x"ca",
    x"5a",
    x"87",
    x"3c",
    x"20",
    x"27",
    x"36",
    x"18",
    x"23",
    x"7e",
    x"c6",
    x"04",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"3d",
    x"fe",
    x"16",
    x"38",
    x"02",
    x"3e",
    x"15",
    x"c6",
    x"60",
    x"77",
    x"3e",
    x"01",
    x"32",
    x"98",
    x"e1",
    x"32",
    x"a0",
    x"e1",
    x"32",
    x"c8",
    x"e1",
    x"21",
    x"2a",
    x"87",
    x"c3",
    x"e3",
    x"86",
    x"3d",
    x"3d",
    x"77",
    x"28",
    x"36",
    x"fe",
    x"10",
    x"28",
    x"07",
    x"fe",
    x"08",
    x"28",
    x"08",
    x"c3",
    x"5a",
    x"87",
    x"21",
    x"3a",
    x"87",
    x"18",
    x"05",
    x"21",
    x"4a",
    x"87",
    x"18",
    x"00",
    x"3a",
    x"17",
    x"e1",
    x"5f",
    x"16",
    x"1a",
    x"06",
    x"04",
    x"c5",
    x"e5",
    x"d5",
    x"01",
    x"04",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"eb",
    x"e1",
    x"0e",
    x"04",
    x"09",
    x"c1",
    x"10",
    x"ea",
    x"c3",
    x"5a",
    x"87",
    x"cd",
    x"0a",
    x"87",
    x"c3",
    x"5a",
    x"87",
    x"3a",
    x"17",
    x"e1",
    x"5f",
    x"16",
    x"1a",
    x"6b",
    x"26",
    x"ef",
    x"06",
    x"04",
    x"c5",
    x"e5",
    x"d5",
    x"01",
    x"04",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"eb",
    x"e1",
    x"09",
    x"c1",
    x"10",
    x"ec",
    x"c9",
    x"c8",
    x"cc",
    x"d2",
    x"ca",
    x"d0",
    x"d4",
    x"d6",
    x"ce",
    x"cd",
    x"d5",
    x"d7",
    x"d3",
    x"c9",
    x"d1",
    x"cf",
    x"cb",
    x"d8",
    x"dc",
    x"e2",
    x"da",
    x"e0",
    x"e4",
    x"e6",
    x"de",
    x"dd",
    x"e5",
    x"e7",
    x"e3",
    x"d9",
    x"e1",
    x"df",
    x"db",
    x"e8",
    x"ec",
    x"f2",
    x"ea",
    x"f0",
    x"f4",
    x"f6",
    x"ee",
    x"ed",
    x"f5",
    x"f7",
    x"f3",
    x"e9",
    x"f1",
    x"ef",
    x"eb",
    x"21",
    x"00",
    x"e1",
    x"11",
    x"e0",
    x"e7",
    x"06",
    x"04",
    x"c5",
    x"e5",
    x"d5",
    x"7e",
    x"a7",
    x"ca",
    x"fd",
    x"87",
    x"fe",
    x"ff",
    x"28",
    x"2e",
    x"3d",
    x"77",
    x"28",
    x"3e",
    x"1c",
    x"1c",
    x"fe",
    x"12",
    x"28",
    x"1b",
    x"fe",
    x"0c",
    x"28",
    x"0e",
    x"fe",
    x"06",
    x"c2",
    x"fd",
    x"87",
    x"3e",
    x"ac",
    x"12",
    x"13",
    x"3e",
    x"0f",
    x"12",
    x"18",
    x"73",
    x"3e",
    x"a8",
    x"12",
    x"13",
    x"3e",
    x"0f",
    x"12",
    x"18",
    x"6a",
    x"3e",
    x"a4",
    x"12",
    x"13",
    x"3e",
    x"0f",
    x"12",
    x"18",
    x"61",
    x"36",
    x"17",
    x"2c",
    x"2c",
    x"7e",
    x"12",
    x"2c",
    x"1c",
    x"7e",
    x"12",
    x"1c",
    x"3e",
    x"a0",
    x"12",
    x"1c",
    x"3e",
    x"0f",
    x"12",
    x"18",
    x"4d",
    x"3e",
    x"e0",
    x"12",
    x"2c",
    x"7e",
    x"36",
    x"00",
    x"fe",
    x"0f",
    x"30",
    x"42",
    x"87",
    x"11",
    x"27",
    x"88",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"a7",
    x"28",
    x"35",
    x"23",
    x"4f",
    x"13",
    x"1a",
    x"47",
    x"e5",
    x"c5",
    x"21",
    x"11",
    x"e1",
    x"11",
    x"f0",
    x"e7",
    x"7e",
    x"3c",
    x"e6",
    x"03",
    x"77",
    x"23",
    x"47",
    x"87",
    x"87",
    x"83",
    x"5f",
    x"78",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"36",
    x"3c",
    x"c1",
    x"e1",
    x"7e",
    x"c6",
    x"04",
    x"fe",
    x"f0",
    x"38",
    x"01",
    x"af",
    x"12",
    x"2c",
    x"1c",
    x"7e",
    x"12",
    x"1c",
    x"79",
    x"12",
    x"1c",
    x"78",
    x"12",
    x"d1",
    x"e1",
    x"7b",
    x"c6",
    x"04",
    x"5f",
    x"7d",
    x"c6",
    x"04",
    x"6f",
    x"c1",
    x"05",
    x"c2",
    x"62",
    x"87",
    x"06",
    x"04",
    x"21",
    x"12",
    x"e1",
    x"11",
    x"f0",
    x"e7",
    x"7e",
    x"a7",
    x"28",
    x"06",
    x"35",
    x"20",
    x"03",
    x"3e",
    x"e0",
    x"12",
    x"2c",
    x"1c",
    x"1c",
    x"1c",
    x"1c",
    x"10",
    x"ef",
    x"18",
    x"1e",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"d4",
    x"0e",
    x"d8",
    x"0b",
    x"e4",
    x"0a",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"dc",
    x"0c",
    x"00",
    x"00",
    x"dc",
    x"07",
    x"e0",
    x"05",
    x"e8",
    x"0d",
    x"ec",
    x"09",
    x"21",
    x"20",
    x"e1",
    x"7e",
    x"a7",
    x"ca",
    x"94",
    x"86",
    x"3a",
    x"b4",
    x"e7",
    x"fe",
    x"e0",
    x"20",
    x"02",
    x"36",
    x"03",
    x"7e",
    x"fe",
    x"02",
    x"28",
    x"74",
    x"47",
    x"23",
    x"7e",
    x"23",
    x"d6",
    x"0c",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"4f",
    x"34",
    x"7e",
    x"23",
    x"be",
    x"da",
    x"94",
    x"86",
    x"2b",
    x"36",
    x"00",
    x"23",
    x"23",
    x"78",
    x"3d",
    x"28",
    x"23",
    x"7e",
    x"a7",
    x"20",
    x"08",
    x"32",
    x"20",
    x"e1",
    x"32",
    x"b8",
    x"e1",
    x"18",
    x"01",
    x"35",
    x"0f",
    x"0f",
    x"0f",
    x"81",
    x"21",
    x"e0",
    x"19",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"eb",
    x"01",
    x"06",
    x"00",
    x"cd",
    x"96",
    x"8a",
    x"c3",
    x"94",
    x"86",
    x"7e",
    x"47",
    x"fe",
    x"06",
    x"38",
    x"07",
    x"3e",
    x"02",
    x"32",
    x"20",
    x"e1",
    x"18",
    x"01",
    x"34",
    x"78",
    x"0f",
    x"0f",
    x"0f",
    x"81",
    x"21",
    x"e0",
    x"19",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"78",
    x"11",
    x"c8",
    x"88",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"06",
    x"06",
    x"cd",
    x"cf",
    x"80",
    x"c3",
    x"94",
    x"86",
    x"98",
    x"90",
    x"96",
    x"9c",
    x"a2",
    x"a8",
    x"ae",
    x"23",
    x"23",
    x"34",
    x"7e",
    x"fe",
    x"78",
    x"da",
    x"94",
    x"86",
    x"36",
    x"00",
    x"2b",
    x"2b",
    x"36",
    x"03",
    x"c3",
    x"94",
    x"86",
    x"cd",
    x"f3",
    x"89",
    x"21",
    x"1b",
    x"46",
    x"06",
    x"03",
    x"c5",
    x"cd",
    x"7e",
    x"8a",
    x"c1",
    x"10",
    x"f9",
    x"cd",
    x"fa",
    x"80",
    x"c9",
    x"3e",
    x"04",
    x"32",
    x"60",
    x"e0",
    x"cd",
    x"90",
    x"97",
    x"cd",
    x"9c",
    x"8a",
    x"cd",
    x"25",
    x"8a",
    x"21",
    x"45",
    x"18",
    x"cd",
    x"46",
    x"86",
    x"21",
    x"52",
    x"18",
    x"cd",
    x"3e",
    x"86",
    x"21",
    x"1b",
    x"89",
    x"06",
    x"0a",
    x"c5",
    x"cd",
    x"7e",
    x"8a",
    x"c1",
    x"10",
    x"f9",
    x"c9",
    x"26",
    x"18",
    x"05",
    x"13",
    x"03",
    x"0f",
    x"12",
    x"05",
    x"31",
    x"18",
    x"08",
    x"08",
    x"09",
    x"1b",
    x"13",
    x"03",
    x"0f",
    x"12",
    x"05",
    x"68",
    x"19",
    x"0e",
    x"80",
    x"85",
    x"83",
    x"78",
    x"25",
    x"83",
    x"80",
    x"71",
    x"73",
    x"75",
    x"00",
    x"7b",
    x"75",
    x"89",
    x"eb",
    x"19",
    x"08",
    x"28",
    x"29",
    x"2a",
    x"2b",
    x"2c",
    x"2d",
    x"2e",
    x"2f",
    x"64",
    x"1a",
    x"16",
    x"5f",
    x"00",
    x"31",
    x"39",
    x"38",
    x"31",
    x"26",
    x"31",
    x"39",
    x"38",
    x"34",
    x"00",
    x"4e",
    x"41",
    x"4d",
    x"43",
    x"4f",
    x"00",
    x"4c",
    x"54",
    x"44",
    x"5d",
    x"a6",
    x"1a",
    x"13",
    x"41",
    x"4c",
    x"4c",
    x"00",
    x"52",
    x"49",
    x"47",
    x"48",
    x"54",
    x"53",
    x"00",
    x"52",
    x"45",
    x"53",
    x"45",
    x"52",
    x"56",
    x"45",
    x"44",
    x"a4",
    x"18",
    x"18",
    x"25",
    x"a1",
    x"a2",
    x"a3",
    x"00",
    x"b1",
    x"b2",
    x"b3",
    x"00",
    x"c1",
    x"25",
    x"23",
    x"00",
    x"b1",
    x"b2",
    x"b3",
    x"25",
    x"a1",
    x"a2",
    x"a3",
    x"00",
    x"b1",
    x"b2",
    x"b3",
    x"c4",
    x"18",
    x"18",
    x"a4",
    x"a5",
    x"a6",
    x"a7",
    x"b4",
    x"b5",
    x"00",
    x"b7",
    x"00",
    x"c5",
    x"26",
    x"20",
    x"b4",
    x"b5",
    x"24",
    x"b7",
    x"a4",
    x"a5",
    x"a6",
    x"a7",
    x"b4",
    x"b5",
    x"00",
    x"b7",
    x"e4",
    x"18",
    x"18",
    x"a8",
    x"a9",
    x"00",
    x"ab",
    x"b8",
    x"b9",
    x"ba",
    x"bb",
    x"00",
    x"c9",
    x"27",
    x"21",
    x"b8",
    x"b9",
    x"ba",
    x"bb",
    x"a8",
    x"a9",
    x"00",
    x"ab",
    x"b8",
    x"b9",
    x"ba",
    x"bb",
    x"04",
    x"19",
    x"18",
    x"00",
    x"ad",
    x"ae",
    x"af",
    x"bc",
    x"bd",
    x"27",
    x"bf",
    x"00",
    x"cd",
    x"ce",
    x"cf",
    x"bc",
    x"bd",
    x"00",
    x"bf",
    x"00",
    x"ad",
    x"ae",
    x"af",
    x"bc",
    x"bd",
    x"27",
    x"bf",
    x"21",
    x"80",
    x"e7",
    x"06",
    x"20",
    x"36",
    x"e0",
    x"7d",
    x"c6",
    x"04",
    x"6f",
    x"10",
    x"f8",
    x"c9",
    x"01",
    x"01",
    x"82",
    x"cd",
    x"47",
    x"00",
    x"21",
    x"00",
    x"18",
    x"01",
    x"00",
    x"03",
    x"af",
    x"cd",
    x"56",
    x"00",
    x"06",
    x"18",
    x"21",
    x"00",
    x"ef",
    x"11",
    x"00",
    x"18",
    x"c5",
    x"d5",
    x"e5",
    x"01",
    x"19",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"7d",
    x"c6",
    x"20",
    x"6f",
    x"d1",
    x"3e",
    x"20",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"c1",
    x"10",
    x"e7",
    x"c9",
    x"06",
    x"18",
    x"21",
    x"00",
    x"ef",
    x"11",
    x"00",
    x"18",
    x"c5",
    x"01",
    x"10",
    x"00",
    x"e5",
    x"d5",
    x"c5",
    x"cd",
    x"5c",
    x"00",
    x"c1",
    x"e1",
    x"09",
    x"eb",
    x"e1",
    x"e5",
    x"d5",
    x"c5",
    x"cd",
    x"5c",
    x"00",
    x"c1",
    x"e1",
    x"09",
    x"eb",
    x"e1",
    x"7d",
    x"c6",
    x"20",
    x"6f",
    x"c1",
    x"10",
    x"df",
    x"c9",
    x"d9",
    x"0e",
    x"60",
    x"18",
    x"03",
    x"d9",
    x"0e",
    x"30",
    x"d9",
    x"1a",
    x"d9",
    x"06",
    x"02",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"f5",
    x"e6",
    x"0f",
    x"d9",
    x"28",
    x"12",
    x"0e",
    x"00",
    x"d9",
    x"81",
    x"d9",
    x"cd",
    x"4d",
    x"00",
    x"23",
    x"d9",
    x"f1",
    x"10",
    x"e9",
    x"d9",
    x"13",
    x"10",
    x"e1",
    x"c9",
    x"0d",
    x"fa",
    x"68",
    x"8a",
    x"18",
    x"ed",
    x"5e",
    x"23",
    x"56",
    x"23",
    x"06",
    x"00",
    x"4e",
    x"23",
    x"e5",
    x"c5",
    x"cd",
    x"5c",
    x"00",
    x"c1",
    x"e1",
    x"09",
    x"c9",
    x"5e",
    x"23",
    x"56",
    x"23",
    x"4e",
    x"06",
    x"00",
    x"6b",
    x"26",
    x"ef",
    x"c3",
    x"5c",
    x"00",
    x"21",
    x"ba",
    x"8a",
    x"18",
    x"03",
    x"21",
    x"b2",
    x"8a",
    x"01",
    x"00",
    x"08",
    x"c5",
    x"46",
    x"cd",
    x"47",
    x"00",
    x"c1",
    x"23",
    x"0c",
    x"10",
    x"f6",
    x"c9",
    x"02",
    x"82",
    x"06",
    x"ff",
    x"03",
    x"36",
    x"07",
    x"00",
    x"00",
    x"82",
    x"06",
    x"70",
    x"00",
    x"36",
    x"07",
    x"00",
    x"d9",
    x"2a",
    x"07",
    x"e0",
    x"7d",
    x"87",
    x"87",
    x"85",
    x"3c",
    x"6f",
    x"7c",
    x"cb",
    x"24",
    x"3e",
    x"00",
    x"47",
    x"17",
    x"cb",
    x"6c",
    x"20",
    x"01",
    x"04",
    x"a8",
    x"84",
    x"67",
    x"ad",
    x"22",
    x"07",
    x"e0",
    x"d9",
    x"c9",
    x"ed",
    x"73",
    x"05",
    x"e0",
    x"f9",
    x"21",
    x"00",
    x"00",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"10",
    x"f6",
    x"ed",
    x"7b",
    x"05",
    x"e0",
    x"c9",
    x"87",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"e9",
    x"af",
    x"11",
    x"10",
    x"27",
    x"ed",
    x"52",
    x"38",
    x"03",
    x"3c",
    x"18",
    x"f9",
    x"19",
    x"eb",
    x"08",
    x"21",
    x"00",
    x"00",
    x"01",
    x"01",
    x"00",
    x"7a",
    x"b3",
    x"28",
    x"18",
    x"cb",
    x"3a",
    x"cb",
    x"1b",
    x"30",
    x"08",
    x"7d",
    x"81",
    x"27",
    x"6f",
    x"7c",
    x"88",
    x"27",
    x"67",
    x"79",
    x"81",
    x"27",
    x"4f",
    x"78",
    x"88",
    x"27",
    x"47",
    x"18",
    x"e4",
    x"08",
    x"eb",
    x"c9",
    x"2a",
    x"f0",
    x"e0",
    x"e5",
    x"cd",
    x"03",
    x"8b",
    x"21",
    x"f6",
    x"e0",
    x"77",
    x"23",
    x"72",
    x"23",
    x"73",
    x"e1",
    x"ed",
    x"5b",
    x"f2",
    x"e0",
    x"af",
    x"ed",
    x"52",
    x"cd",
    x"03",
    x"8b",
    x"21",
    x"f9",
    x"e0",
    x"77",
    x"23",
    x"72",
    x"23",
    x"73",
    x"c9",
    x"11",
    x"fc",
    x"e0",
    x"21",
    x"f8",
    x"e0",
    x"cd",
    x"98",
    x"8b",
    x"a7",
    x"c8",
    x"01",
    x"00",
    x"00",
    x"cd",
    x"a4",
    x"8b",
    x"38",
    x"03",
    x"04",
    x"18",
    x"f8",
    x"cd",
    x"b6",
    x"8b",
    x"13",
    x"cd",
    x"a4",
    x"8b",
    x"38",
    x"03",
    x"0c",
    x"18",
    x"f8",
    x"cd",
    x"8e",
    x"8b",
    x"57",
    x"41",
    x"cd",
    x"8e",
    x"8b",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"21",
    x"fe",
    x"e0",
    x"72",
    x"23",
    x"77",
    x"c9",
    x"78",
    x"a7",
    x"c8",
    x"af",
    x"c6",
    x"01",
    x"27",
    x"10",
    x"fb",
    x"c9",
    x"e5",
    x"c5",
    x"af",
    x"06",
    x"05",
    x"b6",
    x"2b",
    x"10",
    x"fc",
    x"c1",
    x"e1",
    x"c9",
    x"c5",
    x"d5",
    x"e5",
    x"06",
    x"04",
    x"af",
    x"1a",
    x"9e",
    x"27",
    x"12",
    x"1b",
    x"2b",
    x"10",
    x"f8",
    x"e1",
    x"d1",
    x"c1",
    x"c9",
    x"c5",
    x"d5",
    x"e5",
    x"06",
    x"04",
    x"af",
    x"1a",
    x"8e",
    x"27",
    x"12",
    x"1b",
    x"2b",
    x"10",
    x"f8",
    x"e1",
    x"d1",
    x"c1",
    x"c9",
    x"89",
    x"00",
    x"84",
    x"07",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c3",
    x"04",
    x"c5",
    x"2f",
    x"cb",
    x"28",
    x"8c",
    x"cb",
    x"28",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8d",
    x"c4",
    x"50",
    x"82",
    x"d4",
    x"8b",
    x"89",
    x"00",
    x"84",
    x"07",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"82",
    x"06",
    x"8c",
    x"82",
    x"06",
    x"8c",
    x"82",
    x"06",
    x"8c",
    x"88",
    x"01",
    x"82",
    x"f8",
    x"8b",
    x"84",
    x"0b",
    x"38",
    x"c4",
    x"0f",
    x"50",
    x"c9",
    x"25",
    x"58",
    x"c4",
    x"05",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8c",
    x"8d",
    x"83",
    x"89",
    x"00",
    x"84",
    x"07",
    x"88",
    x"01",
    x"c5",
    x"02",
    x"c8",
    x"04",
    x"30",
    x"84",
    x"0b",
    x"68",
    x"85",
    x"10",
    x"84",
    x"01",
    x"8e",
    x"82",
    x"40",
    x"8c",
    x"84",
    x"07",
    x"89",
    x"00",
    x"88",
    x"01",
    x"c5",
    x"02",
    x"c5",
    x"04",
    x"c3",
    x"13",
    x"d7",
    x"04",
    x"3e",
    x"3e",
    x"2a",
    x"2a",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8c",
    x"8d",
    x"82",
    x"51",
    x"8c",
    x"50",
    x"c3",
    x"26",
    x"c3",
    x"05",
    x"82",
    x"38",
    x"8c",
    x"8f",
    x"82",
    x"4a",
    x"8c",
    x"84",
    x"0e",
    x"3f",
    x"89",
    x"00",
    x"88",
    x"01",
    x"c5",
    x"02",
    x"c5",
    x"04",
    x"c3",
    x"13",
    x"d7",
    x"04",
    x"3e",
    x"3e",
    x"2a",
    x"2a",
    x"84",
    x"0b",
    x"c8",
    x"84",
    x"10",
    x"89",
    x"00",
    x"84",
    x"0c",
    x"84",
    x"0e",
    x"10",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"c5",
    x"2f",
    x"cb",
    x"28",
    x"8c",
    x"cb",
    x"28",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8d",
    x"c4",
    x"50",
    x"82",
    x"7c",
    x"8c",
    x"84",
    x"0e",
    x"08",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"c5",
    x"2f",
    x"c2",
    x"28",
    x"48",
    x"84",
    x"05",
    x"89",
    x"00",
    x"84",
    x"0c",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"84",
    x"0b",
    x"54",
    x"c5",
    x"04",
    x"50",
    x"50",
    x"c5",
    x"2f",
    x"cb",
    x"28",
    x"8c",
    x"cb",
    x"28",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8d",
    x"c4",
    x"50",
    x"82",
    x"7c",
    x"8c",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"84",
    x"0b",
    x"54",
    x"c5",
    x"04",
    x"50",
    x"c6",
    x"2f",
    x"50",
    x"84",
    x"05",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"84",
    x"0b",
    x"54",
    x"c5",
    x"04",
    x"82",
    x"dd",
    x"8c",
    x"89",
    x"00",
    x"84",
    x"0c",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"c5",
    x"2f",
    x"cb",
    x"28",
    x"8c",
    x"cb",
    x"28",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8d",
    x"c4",
    x"50",
    x"82",
    x"7c",
    x"8c",
    x"84",
    x"0e",
    x"01",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"2f",
    x"2f",
    x"82",
    x"ee",
    x"5f",
    x"84",
    x"0e",
    x"01",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"2f",
    x"82",
    x"ee",
    x"5f",
    x"86",
    x"78",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c5",
    x"48",
    x"c2",
    x"3f",
    x"cc",
    x"28",
    x"d3",
    x"48",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"c2",
    x"58",
    x"c5",
    x"0d",
    x"58",
    x"58",
    x"cb",
    x"04",
    x"58",
    x"58",
    x"c9",
    x"08",
    x"c3",
    x"50",
    x"84",
    x"05",
    x"86",
    x"50",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c4",
    x"50",
    x"1f",
    x"1f",
    x"85",
    x"1d",
    x"84",
    x"01",
    x"5f",
    x"3f",
    x"30",
    x"c3",
    x"50",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"cb",
    x"48",
    x"d7",
    x"11",
    x"c9",
    x"48",
    x"84",
    x"05",
    x"86",
    x"50",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c4",
    x"50",
    x"c5",
    x"2f",
    x"85",
    x"08",
    x"84",
    x"01",
    x"4f",
    x"c5",
    x"0f",
    x"c8",
    x"48",
    x"84",
    x"05",
    x"86",
    x"50",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c4",
    x"50",
    x"c5",
    x"0f",
    x"85",
    x"18",
    x"84",
    x"01",
    x"4f",
    x"c5",
    x"2f",
    x"c8",
    x"48",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"c3",
    x"50",
    x"85",
    x"18",
    x"84",
    x"01",
    x"c5",
    x"2f",
    x"5f",
    x"cb",
    x"28",
    x"58",
    x"85",
    x"08",
    x"84",
    x"01",
    x"cc",
    x"48",
    x"84",
    x"05",
    x"86",
    x"78",
    x"82",
    x"e2",
    x"8d",
    x"86",
    x"48",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"5f",
    x"85",
    x"18",
    x"84",
    x"01",
    x"cb",
    x"04",
    x"cb",
    x"24",
    x"d7",
    x"04",
    x"cb",
    x"24",
    x"cb",
    x"04",
    x"85",
    x"00",
    x"84",
    x"01",
    x"5f",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"90",
    x"88",
    x"02",
    x"89",
    x"08",
    x"c4",
    x"04",
    x"c5",
    x"50",
    x"c4",
    x"24",
    x"26",
    x"26",
    x"82",
    x"26",
    x"8e",
    x"48",
    x"c3",
    x"2d",
    x"82",
    x"26",
    x"8e",
    x"48",
    x"c3",
    x"2d",
    x"82",
    x"26",
    x"8e",
    x"c6",
    x"24",
    x"c5",
    x"50",
    x"c4",
    x"04",
    x"00",
    x"84",
    x"05",
    x"c3",
    x"26",
    x"58",
    x"cb",
    x"26",
    x"58",
    x"c3",
    x"26",
    x"83",
    x"86",
    x"60",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"48",
    x"c5",
    x"24",
    x"cb",
    x"11",
    x"cb",
    x"0f",
    x"cb",
    x"0d",
    x"cb",
    x"0b",
    x"cb",
    x"08",
    x"cb",
    x"06",
    x"cb",
    x"04",
    x"cb",
    x"02",
    x"84",
    x"0e",
    x"10",
    x"88",
    x"02",
    x"85",
    x"1c",
    x"84",
    x"01",
    x"cc",
    x"48",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"05",
    x"c9",
    x"48",
    x"10",
    x"10",
    x"58",
    x"55",
    x"cf",
    x"06",
    x"58",
    x"0f",
    x"18",
    x"55",
    x"cf",
    x"06",
    x"c6",
    x"4c",
    x"cf",
    x"26",
    x"58",
    x"2f",
    x"30",
    x"10",
    x"18",
    x"5c",
    x"5c",
    x"84",
    x"05",
    x"86",
    x"48",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"50",
    x"82",
    x"94",
    x"8e",
    x"82",
    x"94",
    x"8e",
    x"82",
    x"94",
    x"8e",
    x"5f",
    x"85",
    x"08",
    x"84",
    x"01",
    x"58",
    x"84",
    x"05",
    x"5f",
    x"85",
    x"08",
    x"84",
    x"01",
    x"5f",
    x"85",
    x"10",
    x"84",
    x"01",
    x"83",
    x"86",
    x"08",
    x"87",
    x"90",
    x"88",
    x"02",
    x"89",
    x"06",
    x"c6",
    x"50",
    x"c9",
    x"04",
    x"58",
    x"58",
    x"ca",
    x"24",
    x"5f",
    x"cb",
    x"03",
    x"58",
    x"cb",
    x"22",
    x"50",
    x"85",
    x"00",
    x"84",
    x"01",
    x"50",
    x"84",
    x"05",
    x"86",
    x"48",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"5f",
    x"85",
    x"18",
    x"84",
    x"01",
    x"5f",
    x"85",
    x"0c",
    x"84",
    x"01",
    x"c7",
    x"56",
    x"85",
    x"18",
    x"84",
    x"01",
    x"c8",
    x"51",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"c5",
    x"04",
    x"c5",
    x"50",
    x"c8",
    x"24",
    x"52",
    x"58",
    x"c5",
    x"08",
    x"52",
    x"50",
    x"c8",
    x"24",
    x"c5",
    x"50",
    x"c5",
    x"04",
    x"84",
    x"05",
    x"86",
    x"48",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c7",
    x"4a",
    x"d7",
    x"26",
    x"c2",
    x"16",
    x"d7",
    x"06",
    x"c2",
    x"16",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"58",
    x"c2",
    x"1b",
    x"d7",
    x"08",
    x"5b",
    x"c2",
    x"3b",
    x"84",
    x"05",
    x"f2",
    x"0f",
    x"d1",
    x"78",
    x"88",
    x"98",
    x"b8",
    x"a8",
    x"98",
    x"88",
    x"78",
    x"68",
    x"58",
    x"48",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"08",
    x"18",
    x"28",
    x"38",
    x"48",
    x"38",
    x"28",
    x"18",
    x"08",
    x"b7",
    x"a7",
    x"97",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"28",
    x"48",
    x"68",
    x"78",
    x"98",
    x"b8",
    x"19",
    x"29",
    x"d6",
    x"c0",
    x"d1",
    x"a8",
    x"98",
    x"88",
    x"78",
    x"68",
    x"58",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"38",
    x"48",
    x"58",
    x"c0",
    x"68",
    x"78",
    x"88",
    x"c0",
    x"98",
    x"a8",
    x"b8",
    x"c0",
    x"c0",
    x"c0",
    x"58",
    x"68",
    x"78",
    x"c0",
    x"88",
    x"98",
    x"a8",
    x"c0",
    x"b8",
    x"09",
    x"19",
    x"c0",
    x"c0",
    x"c0",
    x"78",
    x"88",
    x"98",
    x"c0",
    x"a8",
    x"b8",
    x"09",
    x"c0",
    x"19",
    x"29",
    x"39",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"78",
    x"88",
    x"98",
    x"c0",
    x"a8",
    x"b8",
    x"09",
    x"c0",
    x"19",
    x"29",
    x"39",
    x"f5",
    x"f2",
    x"0e",
    x"d2",
    x"78",
    x"48",
    x"68",
    x"28",
    x"48",
    x"08",
    x"28",
    x"b7",
    x"f0",
    x"94",
    x"8f",
    x"f2",
    x"0e",
    x"d1",
    x"08",
    x"38",
    x"68",
    x"98",
    x"09",
    x"98",
    x"68",
    x"38",
    x"f0",
    x"a2",
    x"8f",
    x"f2",
    x"0e",
    x"d4",
    x"48",
    x"28",
    x"48",
    x"78",
    x"b8",
    x"29",
    x"29",
    x"29",
    x"f5",
    x"f2",
    x"0e",
    x"d4",
    x"28",
    x"b7",
    x"28",
    x"48",
    x"78",
    x"b8",
    x"b8",
    x"b8",
    x"f5",
    x"f2",
    x"0e",
    x"d4",
    x"b7",
    x"77",
    x"b7",
    x"28",
    x"48",
    x"68",
    x"68",
    x"68",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"0a",
    x"a9",
    x"f4",
    x"89",
    x"69",
    x"f4",
    x"49",
    x"29",
    x"f4",
    x"09",
    x"a8",
    x"88",
    x"68",
    x"48",
    x"28",
    x"08",
    x"a7",
    x"87",
    x"67",
    x"f4",
    x"47",
    x"27",
    x"f4",
    x"07",
    x"a6",
    x"f5",
    x"f2",
    x"b0",
    x"ee",
    x"c0",
    x"c0",
    x"f5",
    x"f2",
    x"90",
    x"ee",
    x"c0",
    x"c0",
    x"f5",
    x"f2",
    x"50",
    x"d1",
    x"78",
    x"78",
    x"c0",
    x"f0",
    x"fd",
    x"8f",
    x"21",
    x"1a",
    x"90",
    x"18",
    x"03",
    x"21",
    x"1d",
    x"90",
    x"06",
    x"03",
    x"3e",
    x"0b",
    x"f5",
    x"5e",
    x"23",
    x"cd",
    x"93",
    x"00",
    x"f1",
    x"3c",
    x"10",
    x"f6",
    x"c9",
    x"f8",
    x"28",
    x"00",
    x"d4",
    x"06",
    x"00",
    x"21",
    x"80",
    x"e1",
    x"0e",
    x"08",
    x"16",
    x"00",
    x"06",
    x"03",
    x"7a",
    x"5e",
    x"cd",
    x"93",
    x"00",
    x"2c",
    x"3c",
    x"5e",
    x"cd",
    x"93",
    x"00",
    x"2c",
    x"3c",
    x"57",
    x"79",
    x"5e",
    x"cd",
    x"93",
    x"00",
    x"2c",
    x"3c",
    x"4f",
    x"08",
    x"cb",
    x"1e",
    x"cb",
    x"1f",
    x"08",
    x"2c",
    x"10",
    x"e1",
    x"08",
    x"2f",
    x"e6",
    x"e0",
    x"0f",
    x"0f",
    x"f6",
    x"80",
    x"5f",
    x"3e",
    x"07",
    x"cd",
    x"93",
    x"00",
    x"3a",
    x"98",
    x"e1",
    x"3d",
    x"28",
    x"17",
    x"3d",
    x"20",
    x"27",
    x"21",
    x"8d",
    x"e1",
    x"7e",
    x"35",
    x"23",
    x"fe",
    x"ec",
    x"30",
    x"04",
    x"35",
    x"35",
    x"18",
    x"11",
    x"7e",
    x"c6",
    x"08",
    x"77",
    x"18",
    x"0b",
    x"cd",
    x"03",
    x"90",
    x"21",
    x"8d",
    x"e1",
    x"36",
    x"ff",
    x"23",
    x"36",
    x"0a",
    x"5e",
    x"3e",
    x"06",
    x"cd",
    x"93",
    x"00",
    x"18",
    x"07",
    x"3a",
    x"8c",
    x"e1",
    x"a7",
    x"c4",
    x"08",
    x"90",
    x"21",
    x"90",
    x"e1",
    x"06",
    x"01",
    x"cd",
    x"e1",
    x"8a",
    x"21",
    x"90",
    x"e1",
    x"11",
    x"98",
    x"91",
    x"0e",
    x"03",
    x"06",
    x"29",
    x"d5",
    x"e5",
    x"7e",
    x"a7",
    x"c4",
    x"b1",
    x"90",
    x"e1",
    x"11",
    x"08",
    x"00",
    x"19",
    x"d1",
    x"13",
    x"13",
    x"10",
    x"ef",
    x"c9",
    x"3d",
    x"c2",
    x"c4",
    x"90",
    x"e5",
    x"34",
    x"23",
    x"23",
    x"36",
    x"fe",
    x"23",
    x"23",
    x"1a",
    x"77",
    x"13",
    x"23",
    x"1a",
    x"77",
    x"e1",
    x"23",
    x"56",
    x"23",
    x"34",
    x"7e",
    x"ba",
    x"da",
    x"4a",
    x"91",
    x"36",
    x"00",
    x"23",
    x"23",
    x"5e",
    x"23",
    x"56",
    x"1a",
    x"13",
    x"fe",
    x"d0",
    x"da",
    x"3d",
    x"91",
    x"fe",
    x"f0",
    x"38",
    x"31",
    x"e5",
    x"21",
    x"e8",
    x"90",
    x"e6",
    x"0f",
    x"c3",
    x"f8",
    x"8a",
    x"f4",
    x"90",
    x"07",
    x"91",
    x"1b",
    x"91",
    x"25",
    x"91",
    x"2d",
    x"91",
    x"35",
    x"91",
    x"e1",
    x"23",
    x"13",
    x"13",
    x"73",
    x"23",
    x"72",
    x"2b",
    x"2b",
    x"1b",
    x"1a",
    x"1b",
    x"08",
    x"1a",
    x"5f",
    x"08",
    x"57",
    x"18",
    x"cd",
    x"e1",
    x"23",
    x"5e",
    x"23",
    x"56",
    x"2b",
    x"2b",
    x"18",
    x"c4",
    x"e5",
    x"2b",
    x"2b",
    x"2b",
    x"2b",
    x"d6",
    x"d0",
    x"77",
    x"e1",
    x"18",
    x"b9",
    x"e1",
    x"2b",
    x"2b",
    x"1a",
    x"13",
    x"77",
    x"23",
    x"23",
    x"18",
    x"af",
    x"e1",
    x"2b",
    x"2b",
    x"34",
    x"23",
    x"23",
    x"18",
    x"a7",
    x"e1",
    x"2b",
    x"2b",
    x"35",
    x"23",
    x"23",
    x"18",
    x"9f",
    x"e1",
    x"11",
    x"fb",
    x"ff",
    x"19",
    x"36",
    x"00",
    x"c9",
    x"72",
    x"2b",
    x"73",
    x"2b",
    x"7e",
    x"e6",
    x"60",
    x"28",
    x"03",
    x"32",
    x"8c",
    x"e1",
    x"2b",
    x"0d",
    x"f8",
    x"23",
    x"7e",
    x"08",
    x"23",
    x"5e",
    x"23",
    x"56",
    x"1b",
    x"1a",
    x"e6",
    x"f0",
    x"fe",
    x"e0",
    x"28",
    x"38",
    x"21",
    x"ea",
    x"91",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"1a",
    x"e6",
    x"0f",
    x"cb",
    x"3c",
    x"cb",
    x"1d",
    x"3d",
    x"20",
    x"f9",
    x"eb",
    x"79",
    x"87",
    x"87",
    x"21",
    x"80",
    x"e1",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"73",
    x"23",
    x"72",
    x"23",
    x"08",
    x"57",
    x"e6",
    x"1f",
    x"77",
    x"23",
    x"af",
    x"cb",
    x"12",
    x"17",
    x"77",
    x"c9",
    x"21",
    x"00",
    x"00",
    x"18",
    x"df",
    x"d1",
    x"8f",
    x"ee",
    x"8f",
    x"f4",
    x"8f",
    x"ad",
    x"8f",
    x"b9",
    x"8f",
    x"91",
    x"8f",
    x"9f",
    x"8f",
    x"f4",
    x"8f",
    x"02",
    x"92",
    x"30",
    x"95",
    x"1b",
    x"8f",
    x"3e",
    x"8f",
    x"53",
    x"8f",
    x"82",
    x"8f",
    x"a9",
    x"93",
    x"27",
    x"94",
    x"c5",
    x"8f",
    x"14",
    x"92",
    x"4b",
    x"92",
    x"54",
    x"95",
    x"78",
    x"95",
    x"23",
    x"92",
    x"5a",
    x"92",
    x"82",
    x"92",
    x"b8",
    x"92",
    x"fb",
    x"92",
    x"3e",
    x"93",
    x"82",
    x"93",
    x"8f",
    x"93",
    x"9c",
    x"93",
    x"53",
    x"94",
    x"5c",
    x"94",
    x"02",
    x"95",
    x"ba",
    x"94",
    x"b8",
    x"92",
    x"b0",
    x"92",
    x"fa",
    x"8f",
    x"a6",
    x"92",
    x"b5",
    x"93",
    x"e2",
    x"93",
    x"11",
    x"94",
    x"c8",
    x"d5",
    x"c8",
    x"c9",
    x"75",
    x"be",
    x"c4",
    x"b3",
    x"ad",
    x"a9",
    x"28",
    x"a0",
    x"2a",
    x"97",
    x"ae",
    x"8e",
    x"ac",
    x"86",
    x"1d",
    x"7f",
    x"fb",
    x"77",
    x"3f",
    x"71",
    x"f2",
    x"50",
    x"da",
    x"97",
    x"b7",
    x"08",
    x"b7",
    x"97",
    x"87",
    x"67",
    x"87",
    x"97",
    x"57",
    x"47",
    x"07",
    x"97",
    x"97",
    x"f5",
    x"d5",
    x"f0",
    x"38",
    x"92",
    x"96",
    x"b6",
    x"07",
    x"27",
    x"07",
    x"47",
    x"67",
    x"87",
    x"e4",
    x"97",
    x"f5",
    x"d6",
    x"f0",
    x"38",
    x"92",
    x"96",
    x"07",
    x"b6",
    x"27",
    x"07",
    x"47",
    x"27",
    x"57",
    x"47",
    x"97",
    x"87",
    x"97",
    x"b7",
    x"47",
    x"67",
    x"87",
    x"f5",
    x"f2",
    x"50",
    x"48",
    x"08",
    x"28",
    x"b7",
    x"08",
    x"97",
    x"b7",
    x"87",
    x"97",
    x"47",
    x"57",
    x"27",
    x"07",
    x"b6",
    x"96",
    x"86",
    x"f1",
    x"d5",
    x"f0",
    x"6f",
    x"92",
    x"46",
    x"56",
    x"66",
    x"86",
    x"96",
    x"b6",
    x"07",
    x"27",
    x"e4",
    x"47",
    x"f5",
    x"d6",
    x"f0",
    x"6f",
    x"92",
    x"46",
    x"86",
    x"66",
    x"96",
    x"86",
    x"07",
    x"b6",
    x"27",
    x"07",
    x"47",
    x"27",
    x"57",
    x"47",
    x"27",
    x"07",
    x"b6",
    x"f5",
    x"f2",
    x"0d",
    x"08",
    x"97",
    x"b7",
    x"87",
    x"97",
    x"67",
    x"87",
    x"47",
    x"57",
    x"07",
    x"27",
    x"b6",
    x"96",
    x"86",
    x"66",
    x"46",
    x"f1",
    x"d6",
    x"f2",
    x"0d",
    x"95",
    x"95",
    x"46",
    x"46",
    x"96",
    x"96",
    x"96",
    x"46",
    x"26",
    x"06",
    x"b5",
    x"95",
    x"95",
    x"b5",
    x"b5",
    x"b5",
    x"06",
    x"06",
    x"26",
    x"26",
    x"46",
    x"46",
    x"56",
    x"56",
    x"46",
    x"46",
    x"26",
    x"06",
    x"b5",
    x"85",
    x"95",
    x"b5",
    x"f5",
    x"f2",
    x"0b",
    x"d6",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"f0",
    x"bb",
    x"92",
    x"f2",
    x"0d",
    x"d6",
    x"c0",
    x"c0",
    x"f0",
    x"bb",
    x"92",
    x"f2",
    x"0f",
    x"d6",
    x"77",
    x"77",
    x"77",
    x"08",
    x"28",
    x"28",
    x"28",
    x"58",
    x"48",
    x"48",
    x"48",
    x"08",
    x"28",
    x"28",
    x"28",
    x"98",
    x"78",
    x"78",
    x"78",
    x"08",
    x"28",
    x"28",
    x"28",
    x"58",
    x"48",
    x"48",
    x"48",
    x"08",
    x"78",
    x"78",
    x"78",
    x"b8",
    x"09",
    x"09",
    x"09",
    x"a8",
    x"88",
    x"88",
    x"88",
    x"78",
    x"58",
    x"58",
    x"58",
    x"38",
    x"28",
    x"28",
    x"28",
    x"a7",
    x"a8",
    x"a8",
    x"a8",
    x"09",
    x"a8",
    x"a8",
    x"a8",
    x"78",
    x"d8",
    x"98",
    x"58",
    x"28",
    x"78",
    x"48",
    x"28",
    x"f5",
    x"f2",
    x"0d",
    x"d6",
    x"48",
    x"48",
    x"48",
    x"77",
    x"28",
    x"28",
    x"28",
    x"97",
    x"08",
    x"08",
    x"08",
    x"77",
    x"97",
    x"97",
    x"97",
    x"b7",
    x"48",
    x"48",
    x"48",
    x"77",
    x"28",
    x"28",
    x"28",
    x"97",
    x"08",
    x"08",
    x"08",
    x"77",
    x"28",
    x"28",
    x"28",
    x"78",
    x"88",
    x"88",
    x"88",
    x"78",
    x"58",
    x"58",
    x"58",
    x"38",
    x"28",
    x"28",
    x"28",
    x"08",
    x"a7",
    x"a7",
    x"a7",
    x"28",
    x"38",
    x"38",
    x"38",
    x"58",
    x"38",
    x"38",
    x"38",
    x"08",
    x"d8",
    x"58",
    x"28",
    x"97",
    x"28",
    x"b7",
    x"97",
    x"f5",
    x"f2",
    x"0d",
    x"d6",
    x"77",
    x"77",
    x"77",
    x"77",
    x"97",
    x"97",
    x"97",
    x"08",
    x"b7",
    x"b7",
    x"b7",
    x"b7",
    x"77",
    x"77",
    x"77",
    x"77",
    x"08",
    x"08",
    x"08",
    x"08",
    x"28",
    x"28",
    x"28",
    x"58",
    x"48",
    x"48",
    x"48",
    x"48",
    x"28",
    x"28",
    x"28",
    x"28",
    x"38",
    x"38",
    x"38",
    x"38",
    x"28",
    x"28",
    x"28",
    x"08",
    x"a7",
    x"a7",
    x"a7",
    x"a7",
    x"38",
    x"38",
    x"38",
    x"38",
    x"a8",
    x"a8",
    x"a8",
    x"a8",
    x"78",
    x"78",
    x"78",
    x"38",
    x"28",
    x"28",
    x"28",
    x"28",
    x"78",
    x"78",
    x"78",
    x"48",
    x"f5",
    x"f2",
    x"0d",
    x"d7",
    x"28",
    x"28",
    x"c0",
    x"28",
    x"38",
    x"58",
    x"78",
    x"78",
    x"78",
    x"f5",
    x"f2",
    x"0d",
    x"d7",
    x"97",
    x"97",
    x"c0",
    x"97",
    x"a7",
    x"08",
    x"28",
    x"28",
    x"28",
    x"f5",
    x"f2",
    x"0d",
    x"d7",
    x"67",
    x"67",
    x"c0",
    x"67",
    x"77",
    x"97",
    x"b7",
    x"b7",
    x"b7",
    x"f5",
    x"f2",
    x"0f",
    x"d4",
    x"77",
    x"97",
    x"77",
    x"97",
    x"08",
    x"28",
    x"08",
    x"28",
    x"f5",
    x"e8",
    x"f2",
    x"50",
    x"b7",
    x"77",
    x"47",
    x"07",
    x"e2",
    x"c0",
    x"d6",
    x"b7",
    x"e2",
    x"77",
    x"d6",
    x"47",
    x"d8",
    x"07",
    x"47",
    x"77",
    x"37",
    x"67",
    x"97",
    x"e8",
    x"57",
    x"97",
    x"08",
    x"28",
    x"e2",
    x"c0",
    x"d6",
    x"38",
    x"e2",
    x"08",
    x"d6",
    x"87",
    x"d8",
    x"57",
    x"37",
    x"07",
    x"87",
    x"37",
    x"08",
    x"f0",
    x"b5",
    x"93",
    x"e8",
    x"f2",
    x"10",
    x"77",
    x"47",
    x"07",
    x"b6",
    x"d6",
    x"c0",
    x"c0",
    x"c0",
    x"76",
    x"47",
    x"47",
    x"47",
    x"07",
    x"d8",
    x"b6",
    x"07",
    x"47",
    x"07",
    x"37",
    x"57",
    x"e8",
    x"27",
    x"57",
    x"97",
    x"08",
    x"d6",
    x"c0",
    x"c0",
    x"c0",
    x"08",
    x"87",
    x"87",
    x"87",
    x"57",
    x"d8",
    x"37",
    x"07",
    x"86",
    x"57",
    x"37",
    x"86",
    x"f0",
    x"e2",
    x"93",
    x"f2",
    x"0d",
    x"e8",
    x"b7",
    x"b7",
    x"b7",
    x"b7",
    x"b7",
    x"b7",
    x"77",
    x"b7",
    x"97",
    x"97",
    x"97",
    x"97",
    x"87",
    x"87",
    x"08",
    x"28",
    x"f0",
    x"11",
    x"94",
    x"f2",
    x"0e",
    x"d3",
    x"0a",
    x"b9",
    x"a9",
    x"99",
    x"89",
    x"79",
    x"69",
    x"59",
    x"49",
    x"39",
    x"29",
    x"19",
    x"09",
    x"b8",
    x"a8",
    x"98",
    x"88",
    x"78",
    x"68",
    x"58",
    x"48",
    x"38",
    x"28",
    x"18",
    x"08",
    x"b7",
    x"a7",
    x"97",
    x"87",
    x"77",
    x"67",
    x"57",
    x"47",
    x"37",
    x"27",
    x"17",
    x"07",
    x"b6",
    x"a6",
    x"96",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"b8",
    x"c0",
    x"78",
    x"c0",
    x"98",
    x"f5",
    x"d5",
    x"f2",
    x"4f",
    x"48",
    x"48",
    x"f3",
    x"48",
    x"48",
    x"f4",
    x"48",
    x"f3",
    x"48",
    x"f4",
    x"28",
    x"28",
    x"28",
    x"f3",
    x"28",
    x"f4",
    x"28",
    x"28",
    x"28",
    x"f3",
    x"28",
    x"f4",
    x"28",
    x"f3",
    x"28",
    x"d5",
    x"f4",
    x"58",
    x"58",
    x"f3",
    x"58",
    x"58",
    x"f4",
    x"58",
    x"f3",
    x"58",
    x"f4",
    x"48",
    x"48",
    x"48",
    x"f3",
    x"48",
    x"f4",
    x"48",
    x"48",
    x"48",
    x"f3",
    x"48",
    x"f4",
    x"48",
    x"f3",
    x"48",
    x"58",
    x"58",
    x"c0",
    x"58",
    x"f4",
    x"58",
    x"f3",
    x"58",
    x"78",
    x"78",
    x"c0",
    x"78",
    x"f4",
    x"78",
    x"f3",
    x"78",
    x"f4",
    x"78",
    x"f3",
    x"78",
    x"f4",
    x"78",
    x"f3",
    x"78",
    x"98",
    x"98",
    x"c0",
    x"98",
    x"f4",
    x"98",
    x"f3",
    x"98",
    x"f4",
    x"98",
    x"f3",
    x"98",
    x"f0",
    x"27",
    x"94",
    x"f2",
    x"0e",
    x"d5",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"f2",
    x"10",
    x"18",
    x"18",
    x"c0",
    x"18",
    x"f4",
    x"18",
    x"f3",
    x"18",
    x"38",
    x"38",
    x"c0",
    x"38",
    x"f4",
    x"38",
    x"f3",
    x"38",
    x"f4",
    x"38",
    x"f3",
    x"38",
    x"f4",
    x"38",
    x"f3",
    x"38",
    x"f2",
    x"0d",
    x"57",
    x"97",
    x"08",
    x"58",
    x"58",
    x"08",
    x"97",
    x"57",
    x"f5",
    x"f2",
    x"0d",
    x"e4",
    x"07",
    x"76",
    x"07",
    x"76",
    x"07",
    x"76",
    x"07",
    x"76",
    x"d5",
    x"f2",
    x"10",
    x"86",
    x"86",
    x"c0",
    x"86",
    x"f4",
    x"86",
    x"f3",
    x"86",
    x"a6",
    x"a6",
    x"c0",
    x"a6",
    x"f4",
    x"a6",
    x"f3",
    x"a6",
    x"f4",
    x"a6",
    x"f3",
    x"a6",
    x"f4",
    x"a6",
    x"f3",
    x"a6",
    x"f2",
    x"0f",
    x"da",
    x"58",
    x"58",
    x"08",
    x"57",
    x"f5",
    x"f2",
    x"50",
    x"d6",
    x"48",
    x"18",
    x"28",
    x"b7",
    x"08",
    x"97",
    x"b7",
    x"87",
    x"97",
    x"47",
    x"67",
    x"27",
    x"17",
    x"b6",
    x"96",
    x"86",
    x"96",
    x"17",
    x"b6",
    x"27",
    x"17",
    x"47",
    x"27",
    x"67",
    x"47",
    x"97",
    x"87",
    x"97",
    x"b7",
    x"47",
    x"67",
    x"87",
    x"f5",
    x"f2",
    x"0d",
    x"d6",
    x"18",
    x"97",
    x"b7",
    x"87",
    x"97",
    x"67",
    x"87",
    x"47",
    x"67",
    x"17",
    x"27",
    x"b6",
    x"96",
    x"86",
    x"66",
    x"46",
    x"46",
    x"96",
    x"86",
    x"b6",
    x"96",
    x"17",
    x"b6",
    x"27",
    x"17",
    x"47",
    x"27",
    x"67",
    x"47",
    x"27",
    x"17",
    x"b6",
    x"f5",
    x"f2",
    x"0d",
    x"d6",
    x"95",
    x"95",
    x"46",
    x"46",
    x"96",
    x"96",
    x"96",
    x"46",
    x"26",
    x"16",
    x"b5",
    x"95",
    x"95",
    x"b5",
    x"b5",
    x"b5",
    x"16",
    x"16",
    x"26",
    x"26",
    x"46",
    x"46",
    x"66",
    x"66",
    x"46",
    x"46",
    x"26",
    x"16",
    x"b5",
    x"85",
    x"95",
    x"b5",
    x"f5",
    x"fd",
    x"21",
    x"0c",
    x"98",
    x"fd",
    x"7e",
    x"00",
    x"fd",
    x"23",
    x"a7",
    x"ca",
    x"ae",
    x"98",
    x"47",
    x"e6",
    x"3f",
    x"cb",
    x"78",
    x"28",
    x"08",
    x"21",
    x"fd",
    x"95",
    x"cd",
    x"f8",
    x"8a",
    x"18",
    x"e8",
    x"cb",
    x"70",
    x"28",
    x"05",
    x"cd",
    x"17",
    x"96",
    x"18",
    x"df",
    x"cd",
    x"28",
    x"96",
    x"18",
    x"da",
    x"87",
    x"21",
    x"ed",
    x"95",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"7e",
    x"32",
    x"5c",
    x"e0",
    x"23",
    x"e5",
    x"dd",
    x"e1",
    x"11",
    x"00",
    x"f0",
    x"cd",
    x"33",
    x"96",
    x"11",
    x"00",
    x"3c",
    x"21",
    x"00",
    x"f0",
    x"01",
    x"00",
    x"01",
    x"c3",
    x"5c",
    x"00",
    x"4d",
    x"9e",
    x"8f",
    x"9e",
    x"c0",
    x"9e",
    x"f1",
    x"9e",
    x"22",
    x"9f",
    x"64",
    x"9d",
    x"23",
    x"9d",
    x"53",
    x"9f",
    x"33",
    x"96",
    x"80",
    x"96",
    x"b7",
    x"96",
    x"c3",
    x"96",
    x"f0",
    x"96",
    x"d9",
    x"96",
    x"32",
    x"97",
    x"46",
    x"97",
    x"5e",
    x"97",
    x"65",
    x"97",
    x"75",
    x"97",
    x"84",
    x"97",
    x"06",
    x"97",
    x"06",
    x"00",
    x"87",
    x"87",
    x"87",
    x"cb",
    x"10",
    x"4f",
    x"dd",
    x"e5",
    x"e1",
    x"ed",
    x"b0",
    x"e5",
    x"dd",
    x"e1",
    x"c9",
    x"26",
    x"00",
    x"87",
    x"87",
    x"87",
    x"cb",
    x"14",
    x"6f",
    x"19",
    x"eb",
    x"c9",
    x"3e",
    x"02",
    x"cd",
    x"17",
    x"96",
    x"dd",
    x"7e",
    x"00",
    x"3c",
    x"20",
    x"09",
    x"dd",
    x"23",
    x"3e",
    x"06",
    x"cd",
    x"17",
    x"96",
    x"18",
    x"08",
    x"cd",
    x"d9",
    x"96",
    x"3e",
    x"04",
    x"cd",
    x"17",
    x"96",
    x"dd",
    x"7e",
    x"00",
    x"3c",
    x"20",
    x"09",
    x"21",
    x"00",
    x"f0",
    x"01",
    x"c0",
    x"00",
    x"ed",
    x"b0",
    x"c9",
    x"cd",
    x"64",
    x"96",
    x"cd",
    x"64",
    x"96",
    x"cd",
    x"67",
    x"96",
    x"21",
    x"c8",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"d0",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"b0",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"b8",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"c9",
    x"3e",
    x"01",
    x"cd",
    x"17",
    x"96",
    x"21",
    x"08",
    x"00",
    x"19",
    x"d5",
    x"eb",
    x"21",
    x"f0",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"f8",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"d1",
    x"21",
    x"10",
    x"00",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"10",
    x"00",
    x"19",
    x"eb",
    x"c9",
    x"19",
    x"0e",
    x"08",
    x"06",
    x"08",
    x"e5",
    x"cb",
    x"06",
    x"1f",
    x"23",
    x"10",
    x"fa",
    x"e1",
    x"12",
    x"13",
    x"0d",
    x"20",
    x"f1",
    x"c9",
    x"3e",
    x"01",
    x"cd",
    x"28",
    x"96",
    x"3e",
    x"02",
    x"cd",
    x"17",
    x"96",
    x"18",
    x"05",
    x"3e",
    x"03",
    x"cd",
    x"17",
    x"96",
    x"21",
    x"f8",
    x"ff",
    x"cd",
    x"f5",
    x"96",
    x"21",
    x"e8",
    x"ff",
    x"cd",
    x"f5",
    x"96",
    x"21",
    x"d8",
    x"ff",
    x"18",
    x"1c",
    x"21",
    x"f0",
    x"ff",
    x"e5",
    x"cd",
    x"e1",
    x"96",
    x"e1",
    x"cd",
    x"f5",
    x"96",
    x"21",
    x"f8",
    x"ff",
    x"19",
    x"06",
    x"08",
    x"cb",
    x"26",
    x"23",
    x"10",
    x"fb",
    x"c9",
    x"21",
    x"f8",
    x"ff",
    x"18",
    x"ec",
    x"19",
    x"0e",
    x"08",
    x"06",
    x"08",
    x"cb",
    x"06",
    x"1f",
    x"10",
    x"fb",
    x"12",
    x"23",
    x"13",
    x"0d",
    x"20",
    x"f3",
    x"c9",
    x"cd",
    x"12",
    x"97",
    x"cd",
    x"0f",
    x"97",
    x"cd",
    x"0f",
    x"97",
    x"cd",
    x"12",
    x"97",
    x"d5",
    x"21",
    x"d0",
    x"ff",
    x"19",
    x"01",
    x"30",
    x"00",
    x"ed",
    x"b0",
    x"e1",
    x"0e",
    x"06",
    x"af",
    x"08",
    x"af",
    x"06",
    x"08",
    x"08",
    x"cb",
    x"1f",
    x"cb",
    x"1e",
    x"23",
    x"10",
    x"f9",
    x"cb",
    x"1f",
    x"0d",
    x"20",
    x"f1",
    x"c9",
    x"3e",
    x"01",
    x"cd",
    x"17",
    x"96",
    x"3e",
    x"01",
    x"cd",
    x"28",
    x"96",
    x"3e",
    x"01",
    x"cd",
    x"17",
    x"96",
    x"3e",
    x"01",
    x"c3",
    x"28",
    x"96",
    x"3e",
    x"01",
    x"cd",
    x"17",
    x"96",
    x"3e",
    x"01",
    x"cd",
    x"28",
    x"96",
    x"21",
    x"e0",
    x"ff",
    x"19",
    x"01",
    x"08",
    x"00",
    x"ed",
    x"b0",
    x"3e",
    x"01",
    x"c3",
    x"28",
    x"96",
    x"cd",
    x"6a",
    x"97",
    x"e5",
    x"dd",
    x"e1",
    x"c9",
    x"cd",
    x"6a",
    x"97",
    x"eb",
    x"c9",
    x"fd",
    x"6e",
    x"00",
    x"fd",
    x"23",
    x"fd",
    x"66",
    x"00",
    x"fd",
    x"23",
    x"c9",
    x"d5",
    x"cd",
    x"65",
    x"97",
    x"21",
    x"00",
    x"e8",
    x"01",
    x"00",
    x"08",
    x"cd",
    x"5c",
    x"00",
    x"d1",
    x"c9",
    x"21",
    x"00",
    x"f3",
    x"06",
    x"b0",
    x"cd",
    x"e1",
    x"8a",
    x"11",
    x"00",
    x"e8",
    x"c9",
    x"dd",
    x"21",
    x"ec",
    x"97",
    x"11",
    x"00",
    x"f0",
    x"06",
    x"03",
    x"c5",
    x"dd",
    x"6e",
    x"00",
    x"dd",
    x"23",
    x"dd",
    x"66",
    x"00",
    x"dd",
    x"23",
    x"cd",
    x"c2",
    x"97",
    x"c1",
    x"10",
    x"ef",
    x"11",
    x"00",
    x"05",
    x"21",
    x"00",
    x"f0",
    x"01",
    x"80",
    x"01",
    x"cd",
    x"5c",
    x"00",
    x"11",
    x"00",
    x"1c",
    x"21",
    x"f2",
    x"97",
    x"01",
    x"1a",
    x"00",
    x"c3",
    x"5c",
    x"00",
    x"06",
    x"04",
    x"c5",
    x"46",
    x"23",
    x"4e",
    x"23",
    x"3e",
    x"08",
    x"08",
    x"78",
    x"41",
    x"4f",
    x"af",
    x"cb",
    x"11",
    x"30",
    x"02",
    x"f6",
    x"f0",
    x"cb",
    x"11",
    x"30",
    x"02",
    x"f6",
    x"0f",
    x"12",
    x"13",
    x"12",
    x"13",
    x"12",
    x"13",
    x"12",
    x"13",
    x"08",
    x"3d",
    x"20",
    x"e3",
    x"c1",
    x"10",
    x"d9",
    x"c9",
    x"53",
    x"9a",
    x"23",
    x"9a",
    x"7b",
    x"9a",
    x"60",
    x"60",
    x"60",
    x"60",
    x"60",
    x"60",
    x"f0",
    x"f0",
    x"f0",
    x"f0",
    x"f0",
    x"f0",
    x"70",
    x"70",
    x"70",
    x"70",
    x"70",
    x"70",
    x"c0",
    x"40",
    x"40",
    x"40",
    x"40",
    x"40",
    x"40",
    x"40",
    x"8b",
    x"88",
    x"1b",
    x"9a",
    x"60",
    x"08",
    x"88",
    x"7b",
    x"99",
    x"54",
    x"04",
    x"60",
    x"88",
    x"bb",
    x"99",
    x"4c",
    x"04",
    x"60",
    x"88",
    x"d3",
    x"9c",
    x"42",
    x"85",
    x"42",
    x"85",
    x"88",
    x"d3",
    x"9c",
    x"42",
    x"85",
    x"42",
    x"85",
    x"8a",
    x"00",
    x"00",
    x"89",
    x"80",
    x"ec",
    x"88",
    x"1b",
    x"9b",
    x"41",
    x"84",
    x"41",
    x"84",
    x"04",
    x"83",
    x"8a",
    x"00",
    x"08",
    x"89",
    x"80",
    x"ec",
    x"83",
    x"83",
    x"83",
    x"83",
    x"83",
    x"83",
    x"45",
    x"84",
    x"41",
    x"84",
    x"41",
    x"84",
    x"41",
    x"84",
    x"45",
    x"84",
    x"41",
    x"84",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"8a",
    x"00",
    x"10",
    x"8b",
    x"88",
    x"a3",
    x"9c",
    x"80",
    x"88",
    x"e3",
    x"9c",
    x"80",
    x"88",
    x"24",
    x"9d",
    x"80",
    x"88",
    x"65",
    x"9d",
    x"80",
    x"20",
    x"81",
    x"81",
    x"81",
    x"81",
    x"80",
    x"44",
    x"86",
    x"87",
    x"87",
    x"87",
    x"87",
    x"86",
    x"87",
    x"8a",
    x"00",
    x"38",
    x"8b",
    x"89",
    x"00",
    x"e9",
    x"88",
    x"24",
    x"9d",
    x"42",
    x"85",
    x"02",
    x"8c",
    x"89",
    x"80",
    x"ea",
    x"88",
    x"13",
    x"9d",
    x"42",
    x"85",
    x"02",
    x"8c",
    x"89",
    x"00",
    x"ec",
    x"88",
    x"65",
    x"9d",
    x"42",
    x"85",
    x"02",
    x"8c",
    x"89",
    x"80",
    x"ed",
    x"88",
    x"54",
    x"9d",
    x"42",
    x"85",
    x"02",
    x"8c",
    x"00",
    x"11",
    x"e6",
    x"98",
    x"21",
    x"00",
    x"20",
    x"1a",
    x"13",
    x"a7",
    x"c8",
    x"47",
    x"cb",
    x"7f",
    x"28",
    x"10",
    x"e6",
    x"70",
    x"c6",
    x"10",
    x"e5",
    x"6f",
    x"26",
    x"00",
    x"78",
    x"29",
    x"29",
    x"44",
    x"4d",
    x"e1",
    x"18",
    x"0b",
    x"e6",
    x"70",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"3c",
    x"4f",
    x"78",
    x"06",
    x"00",
    x"e6",
    x"0f",
    x"07",
    x"07",
    x"07",
    x"07",
    x"c5",
    x"cd",
    x"56",
    x"00",
    x"c1",
    x"09",
    x"18",
    x"ce",
    x"d6",
    x"df",
    x"d7",
    x"84",
    x"8c",
    x"d9",
    x"d9",
    x"ba",
    x"96",
    x"df",
    x"d7",
    x"8f",
    x"76",
    x"57",
    x"66",
    x"27",
    x"46",
    x"27",
    x"57",
    x"16",
    x"76",
    x"76",
    x"76",
    x"d5",
    x"d5",
    x"ba",
    x"96",
    x"df",
    x"da",
    x"7f",
    x"34",
    x"17",
    x"36",
    x"24",
    x"27",
    x"16",
    x"24",
    x"27",
    x"34",
    x"17",
    x"16",
    x"7f",
    x"76",
    x"06",
    x"24",
    x"27",
    x"36",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"06",
    x"24",
    x"27",
    x"06",
    x"7f",
    x"24",
    x"27",
    x"26",
    x"24",
    x"27",
    x"36",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"06",
    x"24",
    x"27",
    x"06",
    x"24",
    x"27",
    x"16",
    x"24",
    x"17",
    x"36",
    x"24",
    x"27",
    x"36",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"06",
    x"24",
    x"27",
    x"06",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"36",
    x"24",
    x"27",
    x"36",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"06",
    x"24",
    x"27",
    x"06",
    x"24",
    x"27",
    x"16",
    x"24",
    x"47",
    x"06",
    x"24",
    x"37",
    x"26",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"16",
    x"14",
    x"37",
    x"24",
    x"47",
    x"7b",
    x"7b",
    x"79",
    x"79",
    x"74",
    x"74",
    x"74",
    x"74",
    x"7d",
    x"7d",
    x"7d",
    x"7d",
    x"7a",
    x"7a",
    x"7a",
    x"7a",
    x"7c",
    x"7c",
    x"7c",
    x"7c",
    x"ef",
    x"00",
    x"3f",
    x"3f",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"8f",
    x"cf",
    x"c0",
    x"cf",
    x"df",
    x"d8",
    x"df",
    x"cf",
    x"cf",
    x"ef",
    x"6c",
    x"ec",
    x"ec",
    x"6c",
    x"ec",
    x"ec",
    x"f8",
    x"fd",
    x"cd",
    x"cd",
    x"cd",
    x"cd",
    x"cd",
    x"cc",
    x"fe",
    x"fe",
    x"80",
    x"80",
    x"80",
    x"80",
    x"fe",
    x"fe",
    x"7e",
    x"ff",
    x"c3",
    x"c3",
    x"c3",
    x"c3",
    x"ff",
    x"7e",
    x"7f",
    x"7f",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"80",
    x"80",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"1c",
    x"26",
    x"63",
    x"63",
    x"63",
    x"32",
    x"1c",
    x"00",
    x"0c",
    x"1c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"3f",
    x"00",
    x"3e",
    x"63",
    x"07",
    x"1e",
    x"3c",
    x"70",
    x"7f",
    x"00",
    x"3f",
    x"06",
    x"0c",
    x"1e",
    x"03",
    x"63",
    x"3e",
    x"00",
    x"0e",
    x"1e",
    x"36",
    x"66",
    x"7f",
    x"06",
    x"06",
    x"00",
    x"7e",
    x"60",
    x"7e",
    x"03",
    x"03",
    x"63",
    x"3e",
    x"00",
    x"1c",
    x"30",
    x"60",
    x"7e",
    x"61",
    x"61",
    x"3e",
    x"00",
    x"7f",
    x"63",
    x"06",
    x"0c",
    x"18",
    x"18",
    x"18",
    x"00",
    x"3c",
    x"62",
    x"72",
    x"3c",
    x"4f",
    x"43",
    x"3e",
    x"00",
    x"3e",
    x"63",
    x"63",
    x"3f",
    x"03",
    x"06",
    x"3c",
    x"00",
    x"60",
    x"78",
    x"7e",
    x"78",
    x"60",
    x"60",
    x"60",
    x"00",
    x"21",
    x"52",
    x"24",
    x"08",
    x"12",
    x"25",
    x"42",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"1c",
    x"36",
    x"63",
    x"63",
    x"7f",
    x"63",
    x"63",
    x"00",
    x"7e",
    x"63",
    x"63",
    x"7e",
    x"63",
    x"63",
    x"7e",
    x"00",
    x"1e",
    x"33",
    x"60",
    x"60",
    x"60",
    x"33",
    x"1e",
    x"00",
    x"7c",
    x"66",
    x"63",
    x"63",
    x"63",
    x"66",
    x"7c",
    x"00",
    x"3f",
    x"30",
    x"30",
    x"3e",
    x"30",
    x"30",
    x"3f",
    x"00",
    x"7f",
    x"60",
    x"60",
    x"7e",
    x"60",
    x"60",
    x"60",
    x"00",
    x"1f",
    x"30",
    x"60",
    x"67",
    x"63",
    x"33",
    x"1f",
    x"00",
    x"63",
    x"63",
    x"63",
    x"7f",
    x"63",
    x"63",
    x"63",
    x"00",
    x"3f",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"3f",
    x"00",
    x"03",
    x"03",
    x"03",
    x"03",
    x"03",
    x"63",
    x"3e",
    x"00",
    x"63",
    x"66",
    x"6c",
    x"78",
    x"7c",
    x"6e",
    x"67",
    x"00",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"3f",
    x"00",
    x"63",
    x"77",
    x"7f",
    x"7f",
    x"6b",
    x"63",
    x"63",
    x"00",
    x"63",
    x"73",
    x"7b",
    x"7f",
    x"6f",
    x"67",
    x"63",
    x"00",
    x"3e",
    x"63",
    x"63",
    x"63",
    x"63",
    x"63",
    x"3e",
    x"00",
    x"7e",
    x"63",
    x"63",
    x"63",
    x"7e",
    x"60",
    x"60",
    x"00",
    x"3e",
    x"63",
    x"63",
    x"63",
    x"6f",
    x"66",
    x"3d",
    x"00",
    x"7e",
    x"63",
    x"63",
    x"67",
    x"7c",
    x"6e",
    x"67",
    x"00",
    x"3c",
    x"66",
    x"60",
    x"3e",
    x"03",
    x"63",
    x"3e",
    x"00",
    x"3f",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"00",
    x"63",
    x"63",
    x"63",
    x"63",
    x"63",
    x"63",
    x"3e",
    x"00",
    x"63",
    x"63",
    x"63",
    x"77",
    x"3e",
    x"1c",
    x"08",
    x"00",
    x"63",
    x"63",
    x"6b",
    x"7f",
    x"7f",
    x"77",
    x"63",
    x"00",
    x"63",
    x"77",
    x"3e",
    x"1c",
    x"3e",
    x"77",
    x"63",
    x"00",
    x"33",
    x"33",
    x"33",
    x"1e",
    x"0c",
    x"0c",
    x"0c",
    x"00",
    x"7f",
    x"07",
    x"0e",
    x"1c",
    x"38",
    x"70",
    x"7f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"3c",
    x"3c",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"7f",
    x"7f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"18",
    x"18",
    x"00",
    x"18",
    x"3c",
    x"3c",
    x"18",
    x"18",
    x"00",
    x"18",
    x"00",
    x"3c",
    x"42",
    x"9d",
    x"a1",
    x"a1",
    x"9d",
    x"42",
    x"3c",
    x"01",
    x"01",
    x"01",
    x"03",
    x"03",
    x"13",
    x"13",
    x"17",
    x"9e",
    x"9c",
    x"bd",
    x"ff",
    x"ff",
    x"ef",
    x"cd",
    x"81",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"01",
    x"00",
    x"00",
    x"03",
    x"20",
    x"20",
    x"10",
    x"0c",
    x"03",
    x"c0",
    x"38",
    x"07",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"04",
    x"03",
    x"00",
    x"08",
    x"07",
    x"00",
    x"0e",
    x"e0",
    x"1f",
    x"80",
    x"70",
    x"0f",
    x"00",
    x"f0",
    x"0f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"18",
    x"07",
    x"00",
    x"30",
    x"0e",
    x"01",
    x"70",
    x"e0",
    x"1f",
    x"00",
    x"f0",
    x"0f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"0f",
    x"c0",
    x"3c",
    x"03",
    x"00",
    x"f0",
    x"0f",
    x"e0",
    x"c0",
    x"3f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"c0",
    x"3f",
    x"02",
    x"01",
    x"00",
    x"04",
    x"03",
    x"00",
    x"07",
    x"00",
    x"1f",
    x"c0",
    x"3c",
    x"03",
    x"80",
    x"78",
    x"07",
    x"f0",
    x"80",
    x"7f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"c0",
    x"3f",
    x"08",
    x"07",
    x"00",
    x"10",
    x"0f",
    x"00",
    x"3e",
    x"01",
    x"0f",
    x"80",
    x"78",
    x"07",
    x"00",
    x"f0",
    x"0f",
    x"e0",
    x"80",
    x"7f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"c0",
    x"3f",
    x"70",
    x"0f",
    x"00",
    x"60",
    x"1e",
    x"01",
    x"00",
    x"00",
    x"1f",
    x"00",
    x"f0",
    x"0f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"80",
    x"7f",
    x"00",
    x"c0",
    x"3f",
    x"00",
    x"80",
    x"7f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"fe",
    x"fe",
    x"00",
    x"fe",
    x"fe",
    x"00",
    x"fe",
    x"ba",
    x"d6",
    x"6c",
    x"38",
    x"10",
    x"00",
    x"00",
    x"fe",
    x"00",
    x"7c",
    x"60",
    x"7c",
    x"0c",
    x"7c",
    x"00",
    x"fe",
    x"fe",
    x"ba",
    x"54",
    x"28",
    x"10",
    x"00",
    x"00",
    x"7f",
    x"7e",
    x"7c",
    x"46",
    x"72",
    x"60",
    x"78",
    x"72",
    x"3a",
    x"1a",
    x"0e",
    x"07",
    x"03",
    x"01",
    x"ff",
    x"fe",
    x"fc",
    x"e6",
    x"c2",
    x"98",
    x"bc",
    x"9e",
    x"ce",
    x"67",
    x"30",
    x"1b",
    x"08",
    x"07",
    x"03",
    x"01",
    x"ff",
    x"fc",
    x"dc",
    x"8c",
    x"80",
    x"90",
    x"84",
    x"80",
    x"fe",
    x"7e",
    x"96",
    x"62",
    x"02",
    x"12",
    x"42",
    x"02",
    x"aa",
    x"3c",
    x"3c",
    x"18",
    x"0b",
    x"07",
    x"03",
    x"01",
    x"aa",
    x"78",
    x"78",
    x"30",
    x"a0",
    x"c0",
    x"80",
    x"00",
    x"ff",
    x"ff",
    x"c3",
    x"c3",
    x"ff",
    x"c3",
    x"c3",
    x"ff",
    x"e1",
    x"70",
    x"38",
    x"1c",
    x"0e",
    x"07",
    x"03",
    x"01",
    x"00",
    x"00",
    x"60",
    x"10",
    x"0c",
    x"05",
    x"02",
    x"0c",
    x"00",
    x"11",
    x"67",
    x"0e",
    x"1d",
    x"1b",
    x"1b",
    x"0d",
    x"00",
    x"00",
    x"00",
    x"1b",
    x"3f",
    x"3a",
    x"6a",
    x"77",
    x"be",
    x"dd",
    x"d2",
    x"94",
    x"c9",
    x"a2",
    x"88",
    x"d2",
    x"80",
    x"40",
    x"28",
    x"10",
    x"67",
    x"0f",
    x"1a",
    x"1d",
    x"1e",
    x"c7",
    x"22",
    x"ae",
    x"6d",
    x"2e",
    x"1d",
    x"3a",
    x"1e",
    x"3f",
    x"35",
    x"1a",
    x"b5",
    x"ea",
    x"55",
    x"aa",
    x"a8",
    x"5a",
    x"2d",
    x"da",
    x"22",
    x"49",
    x"25",
    x"4a",
    x"00",
    x"00",
    x"20",
    x"12",
    x"09",
    x"05",
    x"02",
    x"0c",
    x"01",
    x"03",
    x"86",
    x"6d",
    x"2d",
    x"66",
    x"2f",
    x"0d",
    x"08",
    x"08",
    x"24",
    x"40",
    x"1f",
    x"3e",
    x"39",
    x"5f",
    x"d2",
    x"14",
    x"2b",
    x"89",
    x"54",
    x"29",
    x"e4",
    x"12",
    x"01",
    x"01",
    x"01",
    x"03",
    x"03",
    x"13",
    x"13",
    x"17",
    x"9e",
    x"9c",
    x"bd",
    x"ff",
    x"ff",
    x"ef",
    x"cd",
    x"81",
    x"00",
    x"00",
    x"00",
    x"09",
    x"12",
    x"26",
    x"7f",
    x"fe",
    x"1f",
    x"1f",
    x"07",
    x"0b",
    x"13",
    x"00",
    x"00",
    x"00",
    x"00",
    x"02",
    x"04",
    x"18",
    x"38",
    x"70",
    x"e0",
    x"40",
    x"48",
    x"f0",
    x"e0",
    x"c8",
    x"d0",
    x"e0",
    x"c0",
    x"80",
    x"02",
    x"02",
    x"1f",
    x"09",
    x"07",
    x"19",
    x"38",
    x"f8",
    x"75",
    x"32",
    x"32",
    x"38",
    x"18",
    x"0c",
    x"06",
    x"02",
    x"02",
    x"02",
    x"1f",
    x"09",
    x"07",
    x"09",
    x"38",
    x"f8",
    x"7d",
    x"5a",
    x"d2",
    x"b0",
    x"90",
    x"90",
    x"f0",
    x"60",
    x"00",
    x"08",
    x"0e",
    x"3e",
    x"77",
    x"ce",
    x"b9",
    x"f3",
    x"e4",
    x"c0",
    x"01",
    x"00",
    x"00",
    x"01",
    x"03",
    x"03",
    x"20",
    x"34",
    x"6a",
    x"ec",
    x"32",
    x"3f",
    x"0c",
    x"88",
    x"d8",
    x"bc",
    x"3c",
    x"6e",
    x"d8",
    x"d8",
    x"30",
    x"e0",
    x"00",
    x"00",
    x"00",
    x"12",
    x"32",
    x"35",
    x"37",
    x"3f",
    x"0c",
    x"1f",
    x"3e",
    x"3b",
    x"19",
    x"00",
    x"00",
    x"00",
    x"09",
    x"00",
    x"00",
    x"00",
    x"12",
    x"72",
    x"75",
    x"77",
    x"3f",
    x"1c",
    x"3f",
    x"7e",
    x"3b",
    x"08",
    x"00",
    x"00",
    x"00",
    x"00",
    x"06",
    x"0f",
    x"0e",
    x"0c",
    x"7d",
    x"7f",
    x"7d",
    x"3e",
    x"2d",
    x"0f",
    x"07",
    x"01",
    x"03",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"20",
    x"c0",
    x"48",
    x"f0",
    x"d0",
    x"e4",
    x"4e",
    x"fe",
    x"fc",
    x"e0",
    x"e0",
    x"e0",
    x"00",
    x"00",
    x"00",
    x"00",
    x"11",
    x"17",
    x"0d",
    x"07",
    x"0c",
    x"0f",
    x"1a",
    x"3a",
    x"3b",
    x"39",
    x"00",
    x"00",
    x"00",
    x"05",
    x"00",
    x"00",
    x"00",
    x"21",
    x"17",
    x"0d",
    x"07",
    x"0c",
    x"1f",
    x"3a",
    x"7a",
    x"73",
    x"71",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"01",
    x"01",
    x"00",
    x"7d",
    x"ff",
    x"fa",
    x"67",
    x"0d",
    x"0b",
    x"0e",
    x"00",
    x"01",
    x"01",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"d0",
    x"60",
    x"f0",
    x"50",
    x"6e",
    x"c0",
    x"60",
    x"e0",
    x"e0",
    x"e0",
    x"e0",
    x"c0",
    x"00",
    x"06",
    x"2c",
    x"20",
    x"5b",
    x"52",
    x"05",
    x"65",
    x"00",
    x"02",
    x"1d",
    x"25",
    x"56",
    x"49",
    x"1e",
    x"25",
    x"00",
    x"66",
    x"89",
    x"63",
    x"2c",
    x"c5",
    x"ba",
    x"25",
    x"00",
    x"32",
    x"6d",
    x"09",
    x"64",
    x"18",
    x"a3",
    x"94",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"01",
    x"03",
    x"03",
    x"01",
    x"01",
    x"01",
    x"01",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"02",
    x"04",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"10",
    x"e0",
    x"e0",
    x"e0",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"40",
    x"40",
    x"e0",
    x"e0",
    x"40",
    x"40",
    x"40",
    x"40",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"02",
    x"02",
    x"07",
    x"07",
    x"02",
    x"02",
    x"02",
    x"02",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"08",
    x"19",
    x"29",
    x"49",
    x"7d",
    x"09",
    x"08",
    x"00",
    x"c6",
    x"29",
    x"29",
    x"29",
    x"29",
    x"29",
    x"c6",
    x"00",
    x"38",
    x"45",
    x"45",
    x"39",
    x"45",
    x"45",
    x"38",
    x"00",
    x"98",
    x"a5",
    x"a5",
    x"a5",
    x"a5",
    x"a5",
    x"98",
    x"00",
    x"bc",
    x"a1",
    x"a1",
    x"b9",
    x"85",
    x"85",
    x"b8",
    x"00",
    x"98",
    x"a1",
    x"a1",
    x"b9",
    x"a5",
    x"a5",
    x"98",
    x"00",
    x"62",
    x"95",
    x"15",
    x"25",
    x"45",
    x"85",
    x"f2",
    x"00",
    x"22",
    x"55",
    x"55",
    x"55",
    x"55",
    x"55",
    x"22",
    x"00",
    x"f2",
    x"15",
    x"65",
    x"15",
    x"15",
    x"95",
    x"62",
    x"0d",
    x"00",
    x"00",
    x"00",
    x"02",
    x"2a",
    x"39",
    x"1b",
    x"1b",
    x"07",
    x"03",
    x"03",
    x"11",
    x"09",
    x"06",
    x"00",
    x"00",
    x"ff",
    x"00",
    x"00",
    x"00",
    x"80",
    x"a8",
    x"38",
    x"b0",
    x"b0",
    x"e0",
    x"80",
    x"80",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"02",
    x"03",
    x"07",
    x"06",
    x"05",
    x"03",
    x"07",
    x"07",
    x"07",
    x"08",
    x"08",
    x"07",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"80",
    x"20",
    x"50",
    x"e0",
    x"c8",
    x"d8",
    x"bc",
    x"70",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"03",
    x"00",
    x"00",
    x"01",
    x"01",
    x"05",
    x"0d",
    x"03",
    x"1f",
    x"1f",
    x"3f",
    x"33",
    x"21",
    x"21",
    x"01",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"0e",
    x"1f",
    x"2f",
    x"03",
    x"03",
    x"03",
    x"04",
    x"08",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"c8",
    x"50",
    x"20",
    x"d8",
    x"c8",
    x"e0",
    x"f0",
    x"70",
    x"70",
    x"20",
    x"40",
    x"00",
    x"00",
    x"0a",
    x"00",
    x"00",
    x"00",
    x"01",
    x"23",
    x"27",
    x"3f",
    x"2b",
    x"37",
    x"1d",
    x"0d",
    x"05",
    x"01",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"06",
    x"0c",
    x"1c",
    x"17",
    x"13",
    x"1f",
    x"1f",
    x"13",
    x"05",
    x"09",
    x"13",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"e0",
    x"e0",
    x"e0",
    x"e0",
    x"e4",
    x"bc",
    x"98",
    x"f0",
    x"00",
    x"00",
    x"00",
    x"07",
    x"00",
    x"00",
    x"06",
    x"02",
    x"01",
    x"fd",
    x"7f",
    x"1d",
    x"01",
    x"01",
    x"01",
    x"01",
    x"01",
    x"00",
    x"00",
    x"00",
    x"04",
    x"06",
    x"0f",
    x"0f",
    x"07",
    x"07",
    x"03",
    x"00",
    x"01",
    x"02",
    x"04",
    x"08",
    x"10",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"10",
    x"30",
    x"9c",
    x"a8",
    x"c0",
    x"f0",
    x"7c",
    x"7e",
    x"3f",
    x"0c",
    x"00",
    x"00",
    x"00",
    x"00",
    x"04",
    x"06",
    x"0e",
    x"1f",
    x"1c",
    x"19",
    x"1c",
    x"5f",
    x"6f",
    x"67",
    x"71",
    x"7b",
    x"7f",
    x"6f",
    x"67",
    x"03",
    x"03",
    x"00",
    x"04",
    x"0d",
    x"1d",
    x"39",
    x"7d",
    x"f9",
    x"d8",
    x"1f",
    x"1f",
    x"0f",
    x"1f",
    x"3b",
    x"30",
    x"00",
    x"00",
    x"7c",
    x"fc",
    x"fb",
    x"87",
    x"97",
    x"c7",
    x"e7",
    x"fe",
    x"7c",
    x"00",
    x"2e",
    x"fc",
    x"f8",
    x"70",
    x"e0",
    x"c0",
    x"06",
    x"80",
    x"50",
    x"20",
    x"50",
    x"08",
    x"05",
    x"03",
    x"03",
    x"1f",
    x"7f",
    x"7d",
    x"f1",
    x"c3",
    x"03",
    x"03",
    x"02",
    x"ff",
    x"20",
    x"60",
    x"e0",
    x"e0",
    x"c2",
    x"de",
    x"fc",
    x"f8",
    x"30",
    x"90",
    x"f8",
    x"bc",
    x"8c",
    x"00",
    x"00",
    x"00",
    x"80",
    x"50",
    x"20",
    x"50",
    x"08",
    x"06",
    x"7f",
    x"ff",
    x"ff",
    x"3f",
    x"03",
    x"03",
    x"03",
    x"03",
    x"03",
    x"02",
    x"10",
    x"30",
    x"70",
    x"70",
    x"f0",
    x"e0",
    x"e0",
    x"c0",
    x"38",
    x"9e",
    x"fe",
    x"fc",
    x"8c",
    x"00",
    x"00",
    x"00",
    x"ff",
    x"42",
    x"59",
    x"20",
    x"46",
    x"55",
    x"4b",
    x"41",
    x"53",
    x"48",
    x"49",
    x"e4",
    x"e5",
    x"e8",
    x"ec",
    x"ec",
    x"f2",
    x"f9",
    x"00",
    x"00",
    x"07",
    x"0e",
    x"14",
    x"14",
    x"18",
    x"1b",
    x"1c",
    x"1c",
    x"1b",
    x"18",
    x"14",
    x"14",
    x"0e",
    x"07",
    x"00",
    x"00",
    x"f9",
    x"f2",
    x"ec",
    x"ec",
    x"e8",
    x"e5",
    x"e4",
    x"d8",
    x"d9",
    x"dd",
    x"e4",
    x"e4",
    x"ec",
    x"f6",
    x"00",
    x"00",
    x"0a",
    x"14",
    x"1c",
    x"1c",
    x"23",
    x"27",
    x"28",
    x"28",
    x"27",
    x"23",
    x"1c",
    x"1c",
    x"14",
    x"0a",
    x"00",
    x"00",
    x"f6",
    x"ec",
    x"e4",
    x"e4",
    x"dd",
    x"d9",
    x"d8",
    x"c8",
    x"ca",
    x"d0",
    x"d8",
    x"d8",
    x"e4",
    x"f2",
    x"00",
    x"00",
    x"0e",
    x"1c",
    x"28",
    x"28",
    x"30",
    x"36",
    x"38",
    x"38",
    x"36",
    x"30",
    x"28",
    x"28",
    x"1c",
    x"0e",
    x"00",
    x"00",
    x"f2",
    x"e4",
    x"d8",
    x"d8",
    x"d0",
    x"ca",
    x"c8",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"74",
    x"e0",
    x"7e",
    x"a7",
    x"28",
    x"f6",
    x"fe",
    x"ff",
    x"28",
    x"0c",
    x"3d",
    x"77",
    x"20",
    x"ee",
    x"21",
    x"75",
    x"81",
    x"cd",
    x"8f",
    x"8a",
    x"18",
    x"e6",
    x"36",
    x"78",
    x"06",
    x"3c",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"c1",
    x"10",
    x"f9",
    x"cd",
    x"de",
    x"80",
    x"21",
    x"71",
    x"e0",
    x"34",
    x"20",
    x"03",
    x"2b",
    x"34",
    x"23",
    x"4e",
    x"23",
    x"23",
    x"7e",
    x"c6",
    x"01",
    x"27",
    x"77",
    x"2b",
    x"7e",
    x"ce",
    x"00",
    x"27",
    x"77",
    x"79",
    x"3c",
    x"e6",
    x"03",
    x"28",
    x"14",
    x"21",
    x"6d",
    x"81",
    x"cd",
    x"7e",
    x"8a",
    x"21",
    x"8e",
    x"19",
    x"11",
    x"72",
    x"e0",
    x"01",
    x"03",
    x"02",
    x"cd",
    x"4f",
    x"8a",
    x"18",
    x"16",
    x"3e",
    x"01",
    x"32",
    x"68",
    x"e2",
    x"32",
    x"70",
    x"e2",
    x"32",
    x"78",
    x"e2",
    x"21",
    x"75",
    x"81",
    x"cd",
    x"7e",
    x"8a",
    x"3e",
    x"78",
    x"32",
    x"74",
    x"e0",
    x"3a",
    x"71",
    x"e0",
    x"4f",
    x"21",
    x"19",
    x"1a",
    x"06",
    x"06",
    x"11",
    x"55",
    x"81",
    x"78",
    x"3d",
    x"87",
    x"87",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"b9",
    x"38",
    x"07",
    x"28",
    x"05",
    x"10",
    x"ec",
    x"c3",
    x"00",
    x"80",
    x"91",
    x"ed",
    x"44",
    x"4f",
    x"3e",
    x"01",
    x"32",
    x"80",
    x"e2",
    x"13",
    x"1a",
    x"47",
    x"85",
    x"e6",
    x"10",
    x"20",
    x"08",
    x"7d",
    x"e6",
    x"e0",
    x"f6",
    x"19",
    x"c6",
    x"40",
    x"6f",
    x"e5",
    x"cd",
    x"be",
    x"80",
    x"e1",
    x"7d",
    x"80",
    x"6f",
    x"06",
    x"08",
    x"e5",
    x"c5",
    x"cd",
    x"6e",
    x"41",
    x"c1",
    x"10",
    x"f9",
    x"e1",
    x"c3",
    x"76",
    x"80",
    x"cd",
    x"c1",
    x"80",
    x"13",
    x"1a",
    x"c5",
    x"e5",
    x"cd",
    x"cf",
    x"80",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"c1",
    x"c9",
    x"4f",
    x"cd",
    x"4d",
    x"00",
    x"23",
    x"0c",
    x"79",
    x"10",
    x"f8",
    x"c9",
    x"21",
    x"19",
    x"19",
    x"18",
    x"03",
    x"21",
    x"19",
    x"1a",
    x"06",
    x"08",
    x"c5",
    x"01",
    x"06",
    x"00",
    x"af",
    x"cd",
    x"56",
    x"00",
    x"7d",
    x"c6",
    x"20",
    x"6f",
    x"c1",
    x"10",
    x"f1",
    x"c9",
    x"21",
    x"0e",
    x"e0",
    x"34",
    x"20",
    x"01",
    x"35",
    x"cd",
    x"d9",
    x"80",
    x"11",
    x"0e",
    x"e0",
    x"1a",
    x"a7",
    x"c8",
    x"fe",
    x"07",
    x"30",
    x"2b",
    x"21",
    x"39",
    x"19",
    x"47",
    x"c5",
    x"e5",
    x"3e",
    x"90",
    x"06",
    x"02",
    x"cd",
    x"cf",
    x"80",
    x"e1",
    x"e5",
    x"11",
    x"20",
    x"00",
    x"19",
    x"3e",
    x"92",
    x"06",
    x"02",
    x"cd",
    x"cf",
    x"80",
    x"e1",
    x"23",
    x"23",
    x"7d",
    x"f6",
    x"e0",
    x"3c",
    x"20",
    x"04",
    x"11",
    x"5a",
    x"00",
    x"19",
    x"c1",
    x"10",
    x"da",
    x"c9",
    x"21",
    x"7c",
    x"19",
    x"01",
    x"01",
    x"01",
    x"cd",
    x"58",
    x"45",
    x"21",
    x"89",
    x"81",
    x"c3",
    x"7e",
    x"8a",
    x"21",
    x"b4",
    x"e7",
    x"36",
    x"a3",
    x"23",
    x"36",
    x"60",
    x"23",
    x"36",
    x"00",
    x"23",
    x"36",
    x"0f",
    x"21",
    x"0e",
    x"e0",
    x"35",
    x"18",
    x"a5",
    x"01",
    x"01",
    x"b4",
    x"b5",
    x"05",
    x"01",
    x"b6",
    x"b7",
    x"0a",
    x"02",
    x"b8",
    x"ba",
    x"14",
    x"02",
    x"bc",
    x"be",
    x"1e",
    x"02",
    x"c0",
    x"c2",
    x"32",
    x"02",
    x"c4",
    x"c6",
    x"89",
    x"19",
    x"05",
    x"83",
    x"84",
    x"71",
    x"77",
    x"75",
    x"85",
    x"19",
    x"11",
    x"73",
    x"78",
    x"71",
    x"7c",
    x"7c",
    x"75",
    x"7e",
    x"77",
    x"79",
    x"7e",
    x"77",
    x"00",
    x"83",
    x"84",
    x"71",
    x"77",
    x"75",
    x"5a",
    x"19",
    x"04",
    x"13",
    x"08",
    x"09",
    x"10",
    x"cd",
    x"6e",
    x"41",
    x"11",
    x"28",
    x"e0",
    x"1a",
    x"a7",
    x"20",
    x"24",
    x"3a",
    x"b4",
    x"e7",
    x"fe",
    x"a3",
    x"20",
    x"1d",
    x"21",
    x"20",
    x"e1",
    x"7e",
    x"fe",
    x"02",
    x"20",
    x"15",
    x"23",
    x"3a",
    x"b5",
    x"e7",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"fe",
    x"1e",
    x"30",
    x"08",
    x"3e",
    x"02",
    x"12",
    x"3e",
    x"01",
    x"32",
    x"18",
    x"e0",
    x"11",
    x"b8",
    x"e7",
    x"cd",
    x"e4",
    x"81",
    x"28",
    x"09",
    x"af",
    x"32",
    x"30",
    x"e1",
    x"3e",
    x"e0",
    x"32",
    x"b8",
    x"e7",
    x"11",
    x"bc",
    x"e7",
    x"cd",
    x"e4",
    x"81",
    x"ca",
    x"c3",
    x"84",
    x"af",
    x"32",
    x"36",
    x"e1",
    x"3e",
    x"e0",
    x"32",
    x"bc",
    x"e7",
    x"c3",
    x"c3",
    x"84",
    x"1a",
    x"fe",
    x"e0",
    x"c8",
    x"08",
    x"1c",
    x"1a",
    x"1d",
    x"d9",
    x"5f",
    x"08",
    x"57",
    x"3a",
    x"28",
    x"e0",
    x"3d",
    x"28",
    x"05",
    x"01",
    x"07",
    x"00",
    x"18",
    x"03",
    x"01",
    x"0f",
    x"02",
    x"21",
    x"80",
    x"e7",
    x"d9",
    x"01",
    x"00",
    x"0c",
    x"3a",
    x"28",
    x"e0",
    x"d6",
    x"05",
    x"fe",
    x"03",
    x"30",
    x"01",
    x"04",
    x"d9",
    x"7a",
    x"96",
    x"f2",
    x"17",
    x"82",
    x"ed",
    x"44",
    x"fe",
    x"06",
    x"d2",
    x"46",
    x"82",
    x"2c",
    x"7b",
    x"80",
    x"96",
    x"f2",
    x"25",
    x"82",
    x"ed",
    x"44",
    x"2d",
    x"b9",
    x"d2",
    x"46",
    x"82",
    x"7d",
    x"d9",
    x"0c",
    x"d6",
    x"80",
    x"87",
    x"87",
    x"c6",
    x"04",
    x"6f",
    x"26",
    x"e4",
    x"7e",
    x"e6",
    x"7f",
    x"32",
    x"32",
    x"e0",
    x"d6",
    x"03",
    x"fe",
    x"03",
    x"d9",
    x"38",
    x"03",
    x"cd",
    x"52",
    x"82",
    x"2c",
    x"2c",
    x"2c",
    x"2c",
    x"d9",
    x"05",
    x"c2",
    x"0f",
    x"82",
    x"c3",
    x"ac",
    x"83",
    x"d9",
    x"af",
    x"32",
    x"30",
    x"e0",
    x"7d",
    x"c6",
    x"05",
    x"6f",
    x"7e",
    x"32",
    x"31",
    x"e0",
    x"fe",
    x"2d",
    x"38",
    x"05",
    x"3e",
    x"01",
    x"32",
    x"30",
    x"e0",
    x"7d",
    x"d6",
    x"09",
    x"6f",
    x"d5",
    x"e5",
    x"7e",
    x"3d",
    x"ca",
    x"08",
    x"83",
    x"3d",
    x"ca",
    x"b2",
    x"82",
    x"3d",
    x"ca",
    x"39",
    x"83",
    x"3d",
    x"ca",
    x"46",
    x"83",
    x"3e",
    x"06",
    x"21",
    x"a9",
    x"e0",
    x"35",
    x"20",
    x"03",
    x"3a",
    x"aa",
    x"e0",
    x"32",
    x"33",
    x"e0",
    x"3e",
    x"01",
    x"32",
    x"e0",
    x"e1",
    x"3a",
    x"30",
    x"e0",
    x"a7",
    x"c2",
    x"63",
    x"83",
    x"21",
    x"10",
    x"e0",
    x"35",
    x"3a",
    x"31",
    x"e0",
    x"fe",
    x"19",
    x"30",
    x"07",
    x"21",
    x"12",
    x"e0",
    x"35",
    x"c3",
    x"63",
    x"83",
    x"21",
    x"13",
    x"e0",
    x"35",
    x"c3",
    x"63",
    x"83",
    x"d9",
    x"2c",
    x"2c",
    x"2c",
    x"7e",
    x"fe",
    x"04",
    x"28",
    x"0f",
    x"3e",
    x"01",
    x"32",
    x"f8",
    x"e1",
    x"36",
    x"04",
    x"2d",
    x"2d",
    x"2d",
    x"d9",
    x"e1",
    x"d1",
    x"d9",
    x"c9",
    x"3e",
    x"01",
    x"32",
    x"f0",
    x"e1",
    x"3e",
    x"78",
    x"32",
    x"1a",
    x"e0",
    x"2d",
    x"2d",
    x"2d",
    x"d9",
    x"3a",
    x"0d",
    x"e0",
    x"fe",
    x"03",
    x"20",
    x"0d",
    x"21",
    x"a9",
    x"e0",
    x"35",
    x"20",
    x"07",
    x"3e",
    x"ff",
    x"32",
    x"33",
    x"e0",
    x"18",
    x"0c",
    x"e5",
    x"e1",
    x"7d",
    x"c6",
    x"0c",
    x"6f",
    x"7e",
    x"c6",
    x"03",
    x"32",
    x"33",
    x"e0",
    x"e1",
    x"e5",
    x"3a",
    x"32",
    x"e0",
    x"fe",
    x"09",
    x"20",
    x"4e",
    x"3e",
    x"03",
    x"32",
    x"20",
    x"e1",
    x"18",
    x"47",
    x"af",
    x"32",
    x"a5",
    x"e0",
    x"3c",
    x"32",
    x"d0",
    x"e1",
    x"32",
    x"18",
    x"e2",
    x"32",
    x"20",
    x"e2",
    x"21",
    x"28",
    x"e0",
    x"7e",
    x"36",
    x"00",
    x"fe",
    x"05",
    x"20",
    x"04",
    x"21",
    x"d7",
    x"e4",
    x"34",
    x"21",
    x"b0",
    x"e7",
    x"7e",
    x"3c",
    x"20",
    x"04",
    x"2c",
    x"2c",
    x"7e",
    x"a7",
    x"3e",
    x"09",
    x"20",
    x"01",
    x"3d",
    x"32",
    x"33",
    x"e0",
    x"18",
    x"2a",
    x"3c",
    x"32",
    x"e8",
    x"e1",
    x"e1",
    x"e5",
    x"3e",
    x"06",
    x"32",
    x"33",
    x"e0",
    x"18",
    x"09",
    x"3c",
    x"32",
    x"e0",
    x"e1",
    x"3e",
    x"07",
    x"32",
    x"33",
    x"e0",
    x"3a",
    x"30",
    x"e0",
    x"a7",
    x"20",
    x"0e",
    x"7e",
    x"21",
    x"0f",
    x"e0",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"35",
    x"21",
    x"10",
    x"e0",
    x"35",
    x"21",
    x"a0",
    x"e0",
    x"34",
    x"21",
    x"33",
    x"e0",
    x"7e",
    x"fe",
    x"ff",
    x"20",
    x"09",
    x"3a",
    x"aa",
    x"e0",
    x"77",
    x"cd",
    x"98",
    x"85",
    x"3e",
    x"03",
    x"cd",
    x"98",
    x"85",
    x"e1",
    x"d1",
    x"36",
    x"00",
    x"d9",
    x"d5",
    x"11",
    x"d7",
    x"e4",
    x"1a",
    x"3d",
    x"12",
    x"3a",
    x"10",
    x"e1",
    x"5f",
    x"c6",
    x"04",
    x"e6",
    x"0f",
    x"32",
    x"10",
    x"e1",
    x"7b",
    x"11",
    x"00",
    x"e1",
    x"83",
    x"5f",
    x"3e",
    x"ff",
    x"12",
    x"1c",
    x"3a",
    x"33",
    x"e0",
    x"12",
    x"1c",
    x"7e",
    x"12",
    x"2c",
    x"1c",
    x"7e",
    x"12",
    x"2d",
    x"d1",
    x"36",
    x"e0",
    x"c9",
    x"d9",
    x"21",
    x"00",
    x"e3",
    x"7a",
    x"d6",
    x"0f",
    x"f2",
    x"b8",
    x"83",
    x"ed",
    x"44",
    x"fe",
    x"06",
    x"30",
    x"71",
    x"d9",
    x"06",
    x"04",
    x"d9",
    x"7e",
    x"a7",
    x"ca",
    x"28",
    x"84",
    x"e5",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7b",
    x"80",
    x"96",
    x"f2",
    x"d2",
    x"83",
    x"ed",
    x"44",
    x"b9",
    x"30",
    x"52",
    x"7d",
    x"d6",
    x"2d",
    x"6f",
    x"7e",
    x"3d",
    x"28",
    x"40",
    x"32",
    x"f0",
    x"e1",
    x"e5",
    x"21",
    x"10",
    x"e0",
    x"35",
    x"21",
    x"11",
    x"e0",
    x"35",
    x"21",
    x"14",
    x"e0",
    x"35",
    x"d5",
    x"c5",
    x"af",
    x"cd",
    x"98",
    x"85",
    x"c1",
    x"d1",
    x"e1",
    x"36",
    x"00",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"d5",
    x"3a",
    x"10",
    x"e1",
    x"5f",
    x"c6",
    x"04",
    x"e6",
    x"0f",
    x"32",
    x"10",
    x"e1",
    x"7b",
    x"11",
    x"00",
    x"e1",
    x"83",
    x"5f",
    x"3e",
    x"ff",
    x"12",
    x"1c",
    x"1c",
    x"1c",
    x"7e",
    x"12",
    x"1d",
    x"3e",
    x"0f",
    x"12",
    x"d1",
    x"18",
    x"07",
    x"36",
    x"02",
    x"3e",
    x"01",
    x"32",
    x"f8",
    x"e1",
    x"d9",
    x"0c",
    x"d9",
    x"e1",
    x"2c",
    x"d9",
    x"10",
    x"93",
    x"d9",
    x"21",
    x"5f",
    x"e3",
    x"3e",
    x"04",
    x"08",
    x"7a",
    x"96",
    x"f2",
    x"3a",
    x"84",
    x"ed",
    x"44",
    x"fe",
    x"06",
    x"d2",
    x"b6",
    x"84",
    x"e5",
    x"7d",
    x"d6",
    x"5a",
    x"6f",
    x"d9",
    x"06",
    x"0a",
    x"d9",
    x"7e",
    x"a7",
    x"28",
    x"64",
    x"e5",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7b",
    x"80",
    x"96",
    x"f2",
    x"59",
    x"84",
    x"ed",
    x"44",
    x"b9",
    x"30",
    x"53",
    x"d5",
    x"e5",
    x"08",
    x"57",
    x"08",
    x"7a",
    x"11",
    x"12",
    x"e0",
    x"21",
    x"15",
    x"e0",
    x"fe",
    x"03",
    x"30",
    x"0b",
    x"13",
    x"23",
    x"3e",
    x"01",
    x"32",
    x"e0",
    x"e1",
    x"3e",
    x"02",
    x"18",
    x"05",
    x"3e",
    x"01",
    x"32",
    x"e8",
    x"e1",
    x"35",
    x"eb",
    x"35",
    x"c5",
    x"cd",
    x"98",
    x"85",
    x"c1",
    x"21",
    x"10",
    x"e0",
    x"35",
    x"21",
    x"10",
    x"e1",
    x"7e",
    x"5e",
    x"c6",
    x"04",
    x"e6",
    x"0f",
    x"77",
    x"16",
    x"e1",
    x"e1",
    x"3e",
    x"ff",
    x"12",
    x"1c",
    x"af",
    x"12",
    x"1c",
    x"1c",
    x"7e",
    x"12",
    x"1d",
    x"7d",
    x"c6",
    x"2d",
    x"6f",
    x"7e",
    x"12",
    x"d1",
    x"e1",
    x"36",
    x"00",
    x"d9",
    x"0c",
    x"d9",
    x"18",
    x"01",
    x"e1",
    x"2c",
    x"d9",
    x"10",
    x"93",
    x"d9",
    x"e1",
    x"7d",
    x"c6",
    x"0a",
    x"6f",
    x"08",
    x"3d",
    x"c2",
    x"32",
    x"84",
    x"d9",
    x"79",
    x"a7",
    x"c9",
    x"3a",
    x"28",
    x"e0",
    x"3d",
    x"fa",
    x"d9",
    x"84",
    x"28",
    x"07",
    x"fe",
    x"03",
    x"30",
    x"09",
    x"c3",
    x"90",
    x"81",
    x"21",
    x"b0",
    x"e7",
    x"cd",
    x"e2",
    x"84",
    x"21",
    x"b4",
    x"e7",
    x"cd",
    x"e2",
    x"84",
    x"c3",
    x"90",
    x"81",
    x"56",
    x"7a",
    x"fe",
    x"a3",
    x"c0",
    x"e5",
    x"2c",
    x"5e",
    x"21",
    x"80",
    x"e7",
    x"06",
    x"0c",
    x"3a",
    x"28",
    x"e0",
    x"d6",
    x"05",
    x"fe",
    x"03",
    x"30",
    x"01",
    x"04",
    x"7a",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"4f",
    x"7b",
    x"2c",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"81",
    x"38",
    x"04",
    x"fe",
    x"0e",
    x"38",
    x"26",
    x"2c",
    x"2c",
    x"2c",
    x"10",
    x"e6",
    x"21",
    x"c0",
    x"e7",
    x"06",
    x"08",
    x"7a",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"4f",
    x"7b",
    x"2c",
    x"96",
    x"30",
    x"02",
    x"ed",
    x"44",
    x"81",
    x"38",
    x"04",
    x"fe",
    x"08",
    x"38",
    x"23",
    x"2c",
    x"2c",
    x"2c",
    x"10",
    x"e6",
    x"e1",
    x"c9",
    x"af",
    x"32",
    x"32",
    x"e0",
    x"2c",
    x"2c",
    x"36",
    x"04",
    x"2d",
    x"2d",
    x"2d",
    x"7d",
    x"d9",
    x"d6",
    x"80",
    x"87",
    x"87",
    x"c6",
    x"04",
    x"6f",
    x"26",
    x"e4",
    x"d9",
    x"cd",
    x"52",
    x"82",
    x"18",
    x"0d",
    x"2d",
    x"36",
    x"e0",
    x"11",
    x"80",
    x"f9",
    x"19",
    x"36",
    x"00",
    x"21",
    x"92",
    x"e0",
    x"35",
    x"e1",
    x"36",
    x"e0",
    x"11",
    x"28",
    x"e0",
    x"1a",
    x"3d",
    x"20",
    x"16",
    x"12",
    x"7d",
    x"fe",
    x"b0",
    x"ca",
    x"85",
    x"85",
    x"36",
    x"a3",
    x"2c",
    x"4e",
    x"11",
    x"b0",
    x"e7",
    x"3e",
    x"e0",
    x"12",
    x"1c",
    x"1a",
    x"77",
    x"18",
    x"0a",
    x"3e",
    x"01",
    x"32",
    x"17",
    x"e0",
    x"32",
    x"18",
    x"e0",
    x"2c",
    x"4e",
    x"21",
    x"16",
    x"e1",
    x"7e",
    x"a7",
    x"28",
    x"05",
    x"e5",
    x"cd",
    x"0a",
    x"87",
    x"e1",
    x"36",
    x"ff",
    x"23",
    x"71",
    x"c9",
    x"87",
    x"21",
    x"c7",
    x"85",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"56",
    x"23",
    x"5e",
    x"3a",
    x"0b",
    x"e0",
    x"3d",
    x"c8",
    x"3e",
    x"01",
    x"32",
    x"44",
    x"e0",
    x"21",
    x"43",
    x"e0",
    x"7e",
    x"83",
    x"27",
    x"77",
    x"2b",
    x"7e",
    x"8a",
    x"27",
    x"77",
    x"2b",
    x"7e",
    x"ce",
    x"00",
    x"27",
    x"77",
    x"2b",
    x"7e",
    x"ce",
    x"00",
    x"27",
    x"77",
    x"c9",
    x"01",
    x"50",
    x"00",
    x"80",
    x"00",
    x"50",
    x"04",
    x"00",
    x"08",
    x"00",
    x"16",
    x"00",
    x"01",
    x"60",
    x"01",
    x"00",
    x"05",
    x"00",
    x"10",
    x"00",
    x"01",
    x"60",
    x"10",
    x"00",
    x"15",
    x"00",
    x"20",
    x"00",
    x"30",
    x"00",
    x"3a",
    x"44",
    x"e0",
    x"3d",
    x"c0",
    x"32",
    x"44",
    x"e0",
    x"cd",
    x"7b",
    x"86",
    x"cd",
    x"3b",
    x"86",
    x"cd",
    x"43",
    x"86",
    x"3a",
    x"45",
    x"e0",
    x"21",
    x"46",
    x"e0",
    x"be",
    x"c8",
    x"3a",
    x"41",
    x"e0",
    x"21",
    x"47",
    x"e0",
    x"be",
    x"c0",
    x"3a",
    x"45",
    x"e0",
    x"a7",
    x"20",
    x"01",
    x"77",
    x"3c",
    x"fe",
    x"ff",
    x"28",
    x"03",
    x"32",
    x"45",
    x"e0",
    x"3a",
    x"48",
    x"e0",
    x"86",
    x"27",
    x"77",
    x"3e",
    x"01",
    x"32",
    x"a8",
    x"e1",
    x"32",
    x"b0",
    x"e1",
    x"32",
    x"10",
    x"e2",
    x"c3",
    x"f3",
    x"80",
    x"3a",
    x"09",
    x"e0",
    x"47",
    x"e6",
    x"0f",
    x"c0",
    x"21",
    x"2a",
    x"46",
    x"cb",
    x"60",
    x"c2",
    x"7e",
    x"8a",
    x"c3",
    x"8f",
    x"8a",
    x"21",
    x"59",
    x"18",
    x"11",
    x"01",
    x"e0",
    x"18",
    x"06",
    x"21",
    x"b9",
    x"18",
    x"11",
    x"40",
    x"e0",
    x"01",
    x"04",
    x"03",
    x"d5",
    x"13",
    x"cd",
    x"54",
    x"8a",
    x"d1",
    x"1a",
    x"a7",
    x"c8",
    x"fe",
    x"07",
    x"30",
    x"0e",
    x"47",
    x"11",
    x"1f",
    x"00",
    x"19",
    x"3e",
    x"3a",
    x"cd",
    x"4d",
    x"00",
    x"2b",
    x"10",
    x"f8",
    x"c9",
    x"11",
    x"1a",
    x"18",
    x"19",
    x"eb",
    x"21",
    x"75",
    x"86",
    x"01",
    x"06",
    x"00",
    x"c3",
    x"5c",
    x"00",
    x"20",
    x"47",
    x"52",
    x"45",
    x"41",
    x"54",
    x"11",
    x"40",
    x"e0",
    x"21",
    x"01",
    x"e0",
    x"06",
    x"04",
    x"1a",
    x"be",
    x"d8",
    x"20",
    x"05",
    x"1c",
    x"2c",
    x"10",
    x"f7",
    x"c9",
    x"1a",
    x"77",
    x"1c",
    x"2c",
    x"10",
    x"fa",
    x"c9",
    x"cd",
    x"6e",
    x"41",
    x"21",
    x"16",
    x"e1",
    x"7e",
    x"a7",
    x"ca",
    x"5a",
    x"87",
    x"3c",
    x"20",
    x"27",
    x"36",
    x"18",
    x"23",
    x"7e",
    x"c6",
    x"04",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"3d",
    x"fe",
    x"16",
    x"38",
    x"02",
    x"3e",
    x"15",
    x"c6",
    x"60",
    x"77",
    x"3e",
    x"01",
    x"32",
    x"98",
    x"e1",
    x"32",
    x"a0",
    x"e1",
    x"32",
    x"c8",
    x"e1",
    x"21",
    x"2a",
    x"87",
    x"c3",
    x"e3",
    x"86",
    x"3d",
    x"3d",
    x"77",
    x"28",
    x"36",
    x"fe",
    x"10",
    x"28",
    x"07",
    x"fe",
    x"08",
    x"28",
    x"08",
    x"c3",
    x"5a",
    x"87",
    x"21",
    x"3a",
    x"87",
    x"18",
    x"05",
    x"21",
    x"4a",
    x"87",
    x"18",
    x"00",
    x"3a",
    x"17",
    x"e1",
    x"5f",
    x"16",
    x"1a",
    x"06",
    x"04",
    x"c5",
    x"e5",
    x"d5",
    x"01",
    x"04",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"eb",
    x"e1",
    x"0e",
    x"04",
    x"09",
    x"c1",
    x"10",
    x"ea",
    x"c3",
    x"5a",
    x"87",
    x"cd",
    x"0a",
    x"87",
    x"c3",
    x"5a",
    x"87",
    x"3a",
    x"17",
    x"e1",
    x"5f",
    x"16",
    x"1a",
    x"6b",
    x"26",
    x"ef",
    x"06",
    x"04",
    x"c5",
    x"e5",
    x"d5",
    x"01",
    x"04",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"01",
    x"20",
    x"00",
    x"09",
    x"eb",
    x"e1",
    x"09",
    x"c1",
    x"10",
    x"ec",
    x"c9",
    x"c8",
    x"cc",
    x"d2",
    x"ca",
    x"d0",
    x"d4",
    x"d6",
    x"ce",
    x"cd",
    x"d5",
    x"d7",
    x"d3",
    x"c9",
    x"d1",
    x"cf",
    x"cb",
    x"d8",
    x"dc",
    x"e2",
    x"da",
    x"e0",
    x"e4",
    x"e6",
    x"de",
    x"dd",
    x"e5",
    x"e7",
    x"e3",
    x"d9",
    x"e1",
    x"df",
    x"db",
    x"e8",
    x"ec",
    x"f2",
    x"ea",
    x"f0",
    x"f4",
    x"f6",
    x"ee",
    x"ed",
    x"f5",
    x"f7",
    x"f3",
    x"e9",
    x"f1",
    x"ef",
    x"eb",
    x"21",
    x"00",
    x"e1",
    x"11",
    x"e0",
    x"e7",
    x"06",
    x"04",
    x"c5",
    x"e5",
    x"d5",
    x"7e",
    x"a7",
    x"ca",
    x"fd",
    x"87",
    x"fe",
    x"ff",
    x"28",
    x"2e",
    x"3d",
    x"77",
    x"28",
    x"3e",
    x"1c",
    x"1c",
    x"fe",
    x"12",
    x"28",
    x"1b",
    x"fe",
    x"0c",
    x"28",
    x"0e",
    x"fe",
    x"06",
    x"c2",
    x"fd",
    x"87",
    x"3e",
    x"ac",
    x"12",
    x"13",
    x"3e",
    x"0f",
    x"12",
    x"18",
    x"73",
    x"3e",
    x"a8",
    x"12",
    x"13",
    x"3e",
    x"0f",
    x"12",
    x"18",
    x"6a",
    x"3e",
    x"a4",
    x"12",
    x"13",
    x"3e",
    x"0f",
    x"12",
    x"18",
    x"61",
    x"36",
    x"17",
    x"2c",
    x"2c",
    x"7e",
    x"12",
    x"2c",
    x"1c",
    x"7e",
    x"12",
    x"1c",
    x"3e",
    x"a0",
    x"12",
    x"1c",
    x"3e",
    x"0f",
    x"12",
    x"18",
    x"4d",
    x"3e",
    x"e0",
    x"12",
    x"2c",
    x"7e",
    x"36",
    x"00",
    x"fe",
    x"0f",
    x"30",
    x"42",
    x"87",
    x"11",
    x"27",
    x"88",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"a7",
    x"28",
    x"35",
    x"23",
    x"4f",
    x"13",
    x"1a",
    x"47",
    x"e5",
    x"c5",
    x"21",
    x"11",
    x"e1",
    x"11",
    x"f0",
    x"e7",
    x"7e",
    x"3c",
    x"e6",
    x"03",
    x"77",
    x"23",
    x"47",
    x"87",
    x"87",
    x"83",
    x"5f",
    x"78",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"36",
    x"3c",
    x"c1",
    x"e1",
    x"7e",
    x"c6",
    x"04",
    x"fe",
    x"f0",
    x"38",
    x"01",
    x"af",
    x"12",
    x"2c",
    x"1c",
    x"7e",
    x"12",
    x"1c",
    x"79",
    x"12",
    x"1c",
    x"78",
    x"12",
    x"d1",
    x"e1",
    x"7b",
    x"c6",
    x"04",
    x"5f",
    x"7d",
    x"c6",
    x"04",
    x"6f",
    x"c1",
    x"05",
    x"c2",
    x"62",
    x"87",
    x"06",
    x"04",
    x"21",
    x"12",
    x"e1",
    x"11",
    x"f0",
    x"e7",
    x"7e",
    x"a7",
    x"28",
    x"06",
    x"35",
    x"20",
    x"03",
    x"3e",
    x"e0",
    x"12",
    x"2c",
    x"1c",
    x"1c",
    x"1c",
    x"1c",
    x"10",
    x"ef",
    x"18",
    x"1e",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"d4",
    x"0e",
    x"d8",
    x"0b",
    x"e4",
    x"0a",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"dc",
    x"0c",
    x"00",
    x"00",
    x"dc",
    x"07",
    x"e0",
    x"05",
    x"e8",
    x"0d",
    x"ec",
    x"09",
    x"21",
    x"20",
    x"e1",
    x"7e",
    x"a7",
    x"ca",
    x"94",
    x"86",
    x"3a",
    x"b4",
    x"e7",
    x"fe",
    x"e0",
    x"20",
    x"02",
    x"36",
    x"03",
    x"7e",
    x"fe",
    x"02",
    x"28",
    x"74",
    x"47",
    x"23",
    x"7e",
    x"23",
    x"d6",
    x"0c",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"4f",
    x"34",
    x"7e",
    x"23",
    x"be",
    x"da",
    x"94",
    x"86",
    x"2b",
    x"36",
    x"00",
    x"23",
    x"23",
    x"78",
    x"3d",
    x"28",
    x"23",
    x"7e",
    x"a7",
    x"20",
    x"08",
    x"32",
    x"20",
    x"e1",
    x"32",
    x"b8",
    x"e1",
    x"18",
    x"01",
    x"35",
    x"0f",
    x"0f",
    x"0f",
    x"81",
    x"21",
    x"e0",
    x"19",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"eb",
    x"01",
    x"06",
    x"00",
    x"cd",
    x"96",
    x"8a",
    x"c3",
    x"94",
    x"86",
    x"7e",
    x"47",
    x"fe",
    x"06",
    x"38",
    x"07",
    x"3e",
    x"02",
    x"32",
    x"20",
    x"e1",
    x"18",
    x"01",
    x"34",
    x"78",
    x"0f",
    x"0f",
    x"0f",
    x"81",
    x"21",
    x"e0",
    x"19",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"78",
    x"11",
    x"c8",
    x"88",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"1a",
    x"06",
    x"06",
    x"cd",
    x"cf",
    x"80",
    x"c3",
    x"94",
    x"86",
    x"98",
    x"90",
    x"96",
    x"9c",
    x"a2",
    x"a8",
    x"ae",
    x"23",
    x"23",
    x"34",
    x"7e",
    x"fe",
    x"78",
    x"da",
    x"94",
    x"86",
    x"36",
    x"00",
    x"2b",
    x"2b",
    x"36",
    x"03",
    x"c3",
    x"94",
    x"86",
    x"cd",
    x"f3",
    x"89",
    x"21",
    x"1b",
    x"46",
    x"06",
    x"03",
    x"c5",
    x"cd",
    x"7e",
    x"8a",
    x"c1",
    x"10",
    x"f9",
    x"cd",
    x"fa",
    x"80",
    x"c9",
    x"3e",
    x"04",
    x"32",
    x"60",
    x"e0",
    x"cd",
    x"90",
    x"97",
    x"cd",
    x"9c",
    x"8a",
    x"cd",
    x"25",
    x"8a",
    x"21",
    x"45",
    x"18",
    x"cd",
    x"46",
    x"86",
    x"21",
    x"52",
    x"18",
    x"cd",
    x"3e",
    x"86",
    x"21",
    x"1b",
    x"89",
    x"06",
    x"0a",
    x"c5",
    x"cd",
    x"7e",
    x"8a",
    x"c1",
    x"10",
    x"f9",
    x"c9",
    x"26",
    x"18",
    x"05",
    x"13",
    x"03",
    x"0f",
    x"12",
    x"05",
    x"31",
    x"18",
    x"08",
    x"08",
    x"09",
    x"1b",
    x"13",
    x"03",
    x"0f",
    x"12",
    x"05",
    x"68",
    x"19",
    x"0e",
    x"80",
    x"85",
    x"83",
    x"78",
    x"25",
    x"83",
    x"80",
    x"71",
    x"73",
    x"75",
    x"00",
    x"7b",
    x"75",
    x"89",
    x"eb",
    x"19",
    x"08",
    x"28",
    x"29",
    x"2a",
    x"2b",
    x"2c",
    x"2d",
    x"2e",
    x"2f",
    x"64",
    x"1a",
    x"16",
    x"5f",
    x"00",
    x"31",
    x"39",
    x"38",
    x"31",
    x"26",
    x"31",
    x"39",
    x"38",
    x"34",
    x"00",
    x"4e",
    x"41",
    x"4d",
    x"43",
    x"4f",
    x"00",
    x"4c",
    x"54",
    x"44",
    x"5d",
    x"a6",
    x"1a",
    x"13",
    x"41",
    x"4c",
    x"4c",
    x"00",
    x"52",
    x"49",
    x"47",
    x"48",
    x"54",
    x"53",
    x"00",
    x"52",
    x"45",
    x"53",
    x"45",
    x"52",
    x"56",
    x"45",
    x"44",
    x"a4",
    x"18",
    x"18",
    x"25",
    x"a1",
    x"a2",
    x"a3",
    x"00",
    x"b1",
    x"b2",
    x"b3",
    x"00",
    x"c1",
    x"25",
    x"23",
    x"00",
    x"b1",
    x"b2",
    x"b3",
    x"25",
    x"a1",
    x"a2",
    x"a3",
    x"00",
    x"b1",
    x"b2",
    x"b3",
    x"c4",
    x"18",
    x"18",
    x"a4",
    x"a5",
    x"a6",
    x"a7",
    x"b4",
    x"b5",
    x"00",
    x"b7",
    x"00",
    x"c5",
    x"26",
    x"20",
    x"b4",
    x"b5",
    x"24",
    x"b7",
    x"a4",
    x"a5",
    x"a6",
    x"a7",
    x"b4",
    x"b5",
    x"00",
    x"b7",
    x"e4",
    x"18",
    x"18",
    x"a8",
    x"a9",
    x"00",
    x"ab",
    x"b8",
    x"b9",
    x"ba",
    x"bb",
    x"00",
    x"c9",
    x"27",
    x"21",
    x"b8",
    x"b9",
    x"ba",
    x"bb",
    x"a8",
    x"a9",
    x"00",
    x"ab",
    x"b8",
    x"b9",
    x"ba",
    x"bb",
    x"04",
    x"19",
    x"18",
    x"00",
    x"ad",
    x"ae",
    x"af",
    x"bc",
    x"bd",
    x"27",
    x"bf",
    x"00",
    x"cd",
    x"ce",
    x"cf",
    x"bc",
    x"bd",
    x"00",
    x"bf",
    x"00",
    x"ad",
    x"ae",
    x"af",
    x"bc",
    x"bd",
    x"27",
    x"bf",
    x"21",
    x"80",
    x"e7",
    x"06",
    x"20",
    x"36",
    x"e0",
    x"7d",
    x"c6",
    x"04",
    x"6f",
    x"10",
    x"f8",
    x"c9",
    x"01",
    x"01",
    x"82",
    x"cd",
    x"47",
    x"00",
    x"21",
    x"00",
    x"18",
    x"01",
    x"00",
    x"03",
    x"af",
    x"cd",
    x"56",
    x"00",
    x"06",
    x"18",
    x"21",
    x"00",
    x"ef",
    x"11",
    x"00",
    x"18",
    x"c5",
    x"d5",
    x"e5",
    x"01",
    x"19",
    x"00",
    x"cd",
    x"5c",
    x"00",
    x"e1",
    x"7d",
    x"c6",
    x"20",
    x"6f",
    x"d1",
    x"3e",
    x"20",
    x"83",
    x"5f",
    x"30",
    x"01",
    x"14",
    x"c1",
    x"10",
    x"e7",
    x"c9",
    x"06",
    x"18",
    x"21",
    x"00",
    x"ef",
    x"11",
    x"00",
    x"18",
    x"c5",
    x"01",
    x"10",
    x"00",
    x"e5",
    x"d5",
    x"c5",
    x"cd",
    x"5c",
    x"00",
    x"c1",
    x"e1",
    x"09",
    x"eb",
    x"e1",
    x"e5",
    x"d5",
    x"c5",
    x"cd",
    x"5c",
    x"00",
    x"c1",
    x"e1",
    x"09",
    x"eb",
    x"e1",
    x"7d",
    x"c6",
    x"20",
    x"6f",
    x"c1",
    x"10",
    x"df",
    x"c9",
    x"d9",
    x"0e",
    x"60",
    x"18",
    x"03",
    x"d9",
    x"0e",
    x"30",
    x"d9",
    x"1a",
    x"d9",
    x"06",
    x"02",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"f5",
    x"e6",
    x"0f",
    x"d9",
    x"28",
    x"12",
    x"0e",
    x"00",
    x"d9",
    x"81",
    x"d9",
    x"cd",
    x"4d",
    x"00",
    x"23",
    x"d9",
    x"f1",
    x"10",
    x"e9",
    x"d9",
    x"13",
    x"10",
    x"e1",
    x"c9",
    x"0d",
    x"fa",
    x"68",
    x"8a",
    x"18",
    x"ed",
    x"5e",
    x"23",
    x"56",
    x"23",
    x"06",
    x"00",
    x"4e",
    x"23",
    x"e5",
    x"c5",
    x"cd",
    x"5c",
    x"00",
    x"c1",
    x"e1",
    x"09",
    x"c9",
    x"5e",
    x"23",
    x"56",
    x"23",
    x"4e",
    x"06",
    x"00",
    x"6b",
    x"26",
    x"ef",
    x"c3",
    x"5c",
    x"00",
    x"21",
    x"ba",
    x"8a",
    x"18",
    x"03",
    x"21",
    x"b2",
    x"8a",
    x"01",
    x"00",
    x"08",
    x"c5",
    x"46",
    x"cd",
    x"47",
    x"00",
    x"c1",
    x"23",
    x"0c",
    x"10",
    x"f6",
    x"c9",
    x"02",
    x"82",
    x"06",
    x"ff",
    x"03",
    x"36",
    x"07",
    x"00",
    x"00",
    x"82",
    x"06",
    x"70",
    x"00",
    x"36",
    x"07",
    x"00",
    x"d9",
    x"2a",
    x"07",
    x"e0",
    x"7d",
    x"87",
    x"87",
    x"85",
    x"3c",
    x"6f",
    x"7c",
    x"cb",
    x"24",
    x"3e",
    x"00",
    x"47",
    x"17",
    x"cb",
    x"6c",
    x"20",
    x"01",
    x"04",
    x"a8",
    x"84",
    x"67",
    x"ad",
    x"22",
    x"07",
    x"e0",
    x"d9",
    x"c9",
    x"ed",
    x"73",
    x"05",
    x"e0",
    x"f9",
    x"21",
    x"00",
    x"00",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"e5",
    x"10",
    x"f6",
    x"ed",
    x"7b",
    x"05",
    x"e0",
    x"c9",
    x"87",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"e9",
    x"af",
    x"11",
    x"10",
    x"27",
    x"ed",
    x"52",
    x"38",
    x"03",
    x"3c",
    x"18",
    x"f9",
    x"19",
    x"eb",
    x"08",
    x"21",
    x"00",
    x"00",
    x"01",
    x"01",
    x"00",
    x"7a",
    x"b3",
    x"28",
    x"18",
    x"cb",
    x"3a",
    x"cb",
    x"1b",
    x"30",
    x"08",
    x"7d",
    x"81",
    x"27",
    x"6f",
    x"7c",
    x"88",
    x"27",
    x"67",
    x"79",
    x"81",
    x"27",
    x"4f",
    x"78",
    x"88",
    x"27",
    x"47",
    x"18",
    x"e4",
    x"08",
    x"eb",
    x"c9",
    x"2a",
    x"f0",
    x"e0",
    x"e5",
    x"cd",
    x"03",
    x"8b",
    x"21",
    x"f6",
    x"e0",
    x"77",
    x"23",
    x"72",
    x"23",
    x"73",
    x"e1",
    x"ed",
    x"5b",
    x"f2",
    x"e0",
    x"af",
    x"ed",
    x"52",
    x"cd",
    x"03",
    x"8b",
    x"21",
    x"f9",
    x"e0",
    x"77",
    x"23",
    x"72",
    x"23",
    x"73",
    x"c9",
    x"11",
    x"fc",
    x"e0",
    x"21",
    x"f8",
    x"e0",
    x"cd",
    x"98",
    x"8b",
    x"a7",
    x"c8",
    x"01",
    x"00",
    x"00",
    x"cd",
    x"a4",
    x"8b",
    x"38",
    x"03",
    x"04",
    x"18",
    x"f8",
    x"cd",
    x"b6",
    x"8b",
    x"13",
    x"cd",
    x"a4",
    x"8b",
    x"38",
    x"03",
    x"0c",
    x"18",
    x"f8",
    x"cd",
    x"8e",
    x"8b",
    x"57",
    x"41",
    x"cd",
    x"8e",
    x"8b",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"21",
    x"fe",
    x"e0",
    x"72",
    x"23",
    x"77",
    x"c9",
    x"78",
    x"a7",
    x"c8",
    x"af",
    x"c6",
    x"01",
    x"27",
    x"10",
    x"fb",
    x"c9",
    x"e5",
    x"c5",
    x"af",
    x"06",
    x"05",
    x"b6",
    x"2b",
    x"10",
    x"fc",
    x"c1",
    x"e1",
    x"c9",
    x"c5",
    x"d5",
    x"e5",
    x"06",
    x"04",
    x"af",
    x"1a",
    x"9e",
    x"27",
    x"12",
    x"1b",
    x"2b",
    x"10",
    x"f8",
    x"e1",
    x"d1",
    x"c1",
    x"c9",
    x"c5",
    x"d5",
    x"e5",
    x"06",
    x"04",
    x"af",
    x"1a",
    x"8e",
    x"27",
    x"12",
    x"1b",
    x"2b",
    x"10",
    x"f8",
    x"e1",
    x"d1",
    x"c1",
    x"c9",
    x"89",
    x"00",
    x"84",
    x"07",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c3",
    x"04",
    x"c5",
    x"2f",
    x"cb",
    x"28",
    x"8c",
    x"cb",
    x"28",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8d",
    x"c4",
    x"50",
    x"82",
    x"d4",
    x"8b",
    x"89",
    x"00",
    x"84",
    x"07",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"82",
    x"06",
    x"8c",
    x"82",
    x"06",
    x"8c",
    x"82",
    x"06",
    x"8c",
    x"88",
    x"01",
    x"82",
    x"f8",
    x"8b",
    x"84",
    x"0b",
    x"38",
    x"c4",
    x"0f",
    x"50",
    x"c9",
    x"25",
    x"58",
    x"c4",
    x"05",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8c",
    x"8d",
    x"83",
    x"89",
    x"00",
    x"84",
    x"07",
    x"88",
    x"01",
    x"c5",
    x"02",
    x"c8",
    x"04",
    x"30",
    x"84",
    x"0b",
    x"68",
    x"85",
    x"10",
    x"84",
    x"01",
    x"8e",
    x"82",
    x"40",
    x"8c",
    x"84",
    x"07",
    x"89",
    x"00",
    x"88",
    x"01",
    x"c5",
    x"02",
    x"c5",
    x"04",
    x"c3",
    x"13",
    x"d7",
    x"04",
    x"3e",
    x"3e",
    x"2a",
    x"2a",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8c",
    x"8d",
    x"82",
    x"51",
    x"8c",
    x"50",
    x"c3",
    x"26",
    x"c3",
    x"05",
    x"82",
    x"38",
    x"8c",
    x"8f",
    x"82",
    x"4a",
    x"8c",
    x"84",
    x"0e",
    x"3f",
    x"89",
    x"00",
    x"88",
    x"01",
    x"c5",
    x"02",
    x"c5",
    x"04",
    x"c3",
    x"13",
    x"d7",
    x"04",
    x"3e",
    x"3e",
    x"2a",
    x"2a",
    x"84",
    x"0b",
    x"c8",
    x"84",
    x"10",
    x"89",
    x"00",
    x"84",
    x"0c",
    x"84",
    x"0e",
    x"10",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"c5",
    x"2f",
    x"cb",
    x"28",
    x"8c",
    x"cb",
    x"28",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8d",
    x"c4",
    x"50",
    x"82",
    x"7c",
    x"8c",
    x"84",
    x"0e",
    x"08",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"c5",
    x"2f",
    x"c2",
    x"28",
    x"48",
    x"84",
    x"05",
    x"89",
    x"00",
    x"84",
    x"0c",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"84",
    x"0b",
    x"54",
    x"c5",
    x"04",
    x"50",
    x"50",
    x"c5",
    x"2f",
    x"cb",
    x"28",
    x"8c",
    x"cb",
    x"28",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8d",
    x"c4",
    x"50",
    x"82",
    x"7c",
    x"8c",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"84",
    x"0b",
    x"54",
    x"c5",
    x"04",
    x"50",
    x"c6",
    x"2f",
    x"50",
    x"84",
    x"05",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"84",
    x"0b",
    x"54",
    x"c5",
    x"04",
    x"82",
    x"dd",
    x"8c",
    x"89",
    x"00",
    x"84",
    x"0c",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"c5",
    x"2f",
    x"cb",
    x"28",
    x"8c",
    x"cb",
    x"28",
    x"84",
    x"0b",
    x"c8",
    x"8b",
    x"8d",
    x"c4",
    x"50",
    x"82",
    x"7c",
    x"8c",
    x"84",
    x"0e",
    x"01",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"2f",
    x"2f",
    x"82",
    x"ee",
    x"5f",
    x"84",
    x"0e",
    x"01",
    x"85",
    x"04",
    x"84",
    x"01",
    x"88",
    x"01",
    x"ce",
    x"02",
    x"04",
    x"84",
    x"0b",
    x"58",
    x"c4",
    x"04",
    x"2f",
    x"82",
    x"ee",
    x"5f",
    x"86",
    x"78",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c5",
    x"48",
    x"c2",
    x"3f",
    x"cc",
    x"28",
    x"d3",
    x"48",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"c2",
    x"58",
    x"c5",
    x"0d",
    x"58",
    x"58",
    x"cb",
    x"04",
    x"58",
    x"58",
    x"c9",
    x"08",
    x"c3",
    x"50",
    x"84",
    x"05",
    x"86",
    x"50",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c4",
    x"50",
    x"1f",
    x"1f",
    x"85",
    x"1d",
    x"84",
    x"01",
    x"5f",
    x"3f",
    x"30",
    x"c3",
    x"50",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"cb",
    x"48",
    x"d7",
    x"11",
    x"c9",
    x"48",
    x"84",
    x"05",
    x"86",
    x"50",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c4",
    x"50",
    x"c5",
    x"2f",
    x"85",
    x"08",
    x"84",
    x"01",
    x"4f",
    x"c5",
    x"0f",
    x"c8",
    x"48",
    x"84",
    x"05",
    x"86",
    x"50",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c4",
    x"50",
    x"c5",
    x"0f",
    x"85",
    x"18",
    x"84",
    x"01",
    x"4f",
    x"c5",
    x"2f",
    x"c8",
    x"48",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"c3",
    x"50",
    x"85",
    x"18",
    x"84",
    x"01",
    x"c5",
    x"2f",
    x"5f",
    x"cb",
    x"28",
    x"58",
    x"85",
    x"08",
    x"84",
    x"01",
    x"cc",
    x"48",
    x"84",
    x"05",
    x"86",
    x"78",
    x"82",
    x"e2",
    x"8d",
    x"86",
    x"48",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"5f",
    x"85",
    x"18",
    x"84",
    x"01",
    x"cb",
    x"04",
    x"cb",
    x"24",
    x"d7",
    x"04",
    x"cb",
    x"24",
    x"cb",
    x"04",
    x"85",
    x"00",
    x"84",
    x"01",
    x"5f",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"90",
    x"88",
    x"02",
    x"89",
    x"08",
    x"c4",
    x"04",
    x"c5",
    x"50",
    x"c4",
    x"24",
    x"26",
    x"26",
    x"82",
    x"26",
    x"8e",
    x"48",
    x"c3",
    x"2d",
    x"82",
    x"26",
    x"8e",
    x"48",
    x"c3",
    x"2d",
    x"82",
    x"26",
    x"8e",
    x"c6",
    x"24",
    x"c5",
    x"50",
    x"c4",
    x"04",
    x"00",
    x"84",
    x"05",
    x"c3",
    x"26",
    x"58",
    x"cb",
    x"26",
    x"58",
    x"c3",
    x"26",
    x"83",
    x"86",
    x"60",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"48",
    x"c5",
    x"24",
    x"cb",
    x"11",
    x"cb",
    x"0f",
    x"cb",
    x"0d",
    x"cb",
    x"0b",
    x"cb",
    x"08",
    x"cb",
    x"06",
    x"cb",
    x"04",
    x"cb",
    x"02",
    x"84",
    x"0e",
    x"10",
    x"88",
    x"02",
    x"85",
    x"1c",
    x"84",
    x"01",
    x"cc",
    x"48",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"05",
    x"c9",
    x"48",
    x"10",
    x"10",
    x"58",
    x"55",
    x"cf",
    x"06",
    x"58",
    x"0f",
    x"18",
    x"55",
    x"cf",
    x"06",
    x"c6",
    x"4c",
    x"cf",
    x"26",
    x"58",
    x"2f",
    x"30",
    x"10",
    x"18",
    x"5c",
    x"5c",
    x"84",
    x"05",
    x"86",
    x"48",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"50",
    x"82",
    x"94",
    x"8e",
    x"82",
    x"94",
    x"8e",
    x"82",
    x"94",
    x"8e",
    x"5f",
    x"85",
    x"08",
    x"84",
    x"01",
    x"58",
    x"84",
    x"05",
    x"5f",
    x"85",
    x"08",
    x"84",
    x"01",
    x"5f",
    x"85",
    x"10",
    x"84",
    x"01",
    x"83",
    x"86",
    x"08",
    x"87",
    x"90",
    x"88",
    x"02",
    x"89",
    x"06",
    x"c6",
    x"50",
    x"c9",
    x"04",
    x"58",
    x"58",
    x"ca",
    x"24",
    x"5f",
    x"cb",
    x"03",
    x"58",
    x"cb",
    x"22",
    x"50",
    x"85",
    x"00",
    x"84",
    x"01",
    x"50",
    x"84",
    x"05",
    x"86",
    x"48",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"5f",
    x"85",
    x"18",
    x"84",
    x"01",
    x"5f",
    x"85",
    x"0c",
    x"84",
    x"01",
    x"c7",
    x"56",
    x"85",
    x"18",
    x"84",
    x"01",
    x"c8",
    x"51",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"c5",
    x"04",
    x"c5",
    x"50",
    x"c8",
    x"24",
    x"52",
    x"58",
    x"c5",
    x"08",
    x"52",
    x"50",
    x"c8",
    x"24",
    x"c5",
    x"50",
    x"c5",
    x"04",
    x"84",
    x"05",
    x"86",
    x"48",
    x"87",
    x"ef",
    x"88",
    x"02",
    x"89",
    x"10",
    x"c7",
    x"4a",
    x"d7",
    x"26",
    x"c2",
    x"16",
    x"d7",
    x"06",
    x"c2",
    x"16",
    x"84",
    x"05",
    x"86",
    x"08",
    x"87",
    x"88",
    x"88",
    x"02",
    x"89",
    x"08",
    x"58",
    x"c2",
    x"1b",
    x"d7",
    x"08",
    x"5b",
    x"c2",
    x"3b",
    x"84",
    x"05",
    x"f2",
    x"0f",
    x"d1",
    x"78",
    x"88",
    x"98",
    x"b8",
    x"a8",
    x"98",
    x"88",
    x"78",
    x"68",
    x"58",
    x"48",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"08",
    x"18",
    x"28",
    x"38",
    x"48",
    x"38",
    x"28",
    x"18",
    x"08",
    x"b7",
    x"a7",
    x"97",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"28",
    x"48",
    x"68",
    x"78",
    x"98",
    x"b8",
    x"19",
    x"29",
    x"d6",
    x"c0",
    x"d1",
    x"a8",
    x"98",
    x"88",
    x"78",
    x"68",
    x"58",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"38",
    x"48",
    x"58",
    x"c0",
    x"68",
    x"78",
    x"88",
    x"c0",
    x"98",
    x"a8",
    x"b8",
    x"c0",
    x"c0",
    x"c0",
    x"58",
    x"68",
    x"78",
    x"c0",
    x"88",
    x"98",
    x"a8",
    x"c0",
    x"b8",
    x"09",
    x"19",
    x"c0",
    x"c0",
    x"c0",
    x"78",
    x"88",
    x"98",
    x"c0",
    x"a8",
    x"b8",
    x"09",
    x"c0",
    x"19",
    x"29",
    x"39",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"78",
    x"88",
    x"98",
    x"c0",
    x"a8",
    x"b8",
    x"09",
    x"c0",
    x"19",
    x"29",
    x"39",
    x"f5",
    x"f2",
    x"0e",
    x"d2",
    x"78",
    x"48",
    x"68",
    x"28",
    x"48",
    x"08",
    x"28",
    x"b7",
    x"f0",
    x"94",
    x"8f",
    x"f2",
    x"0e",
    x"d1",
    x"08",
    x"38",
    x"68",
    x"98",
    x"09",
    x"98",
    x"68",
    x"38",
    x"f0",
    x"a2",
    x"8f",
    x"f2",
    x"0e",
    x"d4",
    x"48",
    x"28",
    x"48",
    x"78",
    x"b8",
    x"29",
    x"29",
    x"29",
    x"f5",
    x"f2",
    x"0e",
    x"d4",
    x"28",
    x"b7",
    x"28",
    x"48",
    x"78",
    x"b8",
    x"b8",
    x"b8",
    x"f5",
    x"f2",
    x"0e",
    x"d4",
    x"b7",
    x"77",
    x"b7",
    x"28",
    x"48",
    x"68",
    x"68",
    x"68",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"0a",
    x"a9",
    x"f4",
    x"89",
    x"69",
    x"f4",
    x"49",
    x"29",
    x"f4",
    x"09",
    x"a8",
    x"88",
    x"68",
    x"48",
    x"28",
    x"08",
    x"a7",
    x"87",
    x"67",
    x"f4",
    x"47",
    x"27",
    x"f4",
    x"07",
    x"a6",
    x"f5",
    x"f2",
    x"b0",
    x"ee",
    x"c0",
    x"c0",
    x"f5",
    x"f2",
    x"90",
    x"ee",
    x"c0",
    x"c0",
    x"f5",
    x"f2",
    x"50",
    x"d1",
    x"78",
    x"78",
    x"c0",
    x"f0",
    x"fd",
    x"8f",
    x"21",
    x"1a",
    x"90",
    x"18",
    x"03",
    x"21",
    x"1d",
    x"90",
    x"06",
    x"03",
    x"3e",
    x"0b",
    x"f5",
    x"5e",
    x"23",
    x"cd",
    x"93",
    x"00",
    x"f1",
    x"3c",
    x"10",
    x"f6",
    x"c9",
    x"f8",
    x"28",
    x"00",
    x"d4",
    x"06",
    x"00",
    x"21",
    x"80",
    x"e1",
    x"0e",
    x"08",
    x"16",
    x"00",
    x"06",
    x"03",
    x"7a",
    x"5e",
    x"cd",
    x"93",
    x"00",
    x"2c",
    x"3c",
    x"5e",
    x"cd",
    x"93",
    x"00",
    x"2c",
    x"3c",
    x"57",
    x"79",
    x"5e",
    x"cd",
    x"93",
    x"00",
    x"2c",
    x"3c",
    x"4f",
    x"08",
    x"cb",
    x"1e",
    x"cb",
    x"1f",
    x"08",
    x"2c",
    x"10",
    x"e1",
    x"08",
    x"2f",
    x"e6",
    x"e0",
    x"0f",
    x"0f",
    x"f6",
    x"80",
    x"5f",
    x"3e",
    x"07",
    x"cd",
    x"93",
    x"00",
    x"3a",
    x"98",
    x"e1",
    x"3d",
    x"28",
    x"17",
    x"3d",
    x"20",
    x"27",
    x"21",
    x"8d",
    x"e1",
    x"7e",
    x"35",
    x"23",
    x"fe",
    x"ec",
    x"30",
    x"04",
    x"35",
    x"35",
    x"18",
    x"11",
    x"7e",
    x"c6",
    x"08",
    x"77",
    x"18",
    x"0b",
    x"cd",
    x"03",
    x"90",
    x"21",
    x"8d",
    x"e1",
    x"36",
    x"ff",
    x"23",
    x"36",
    x"0a",
    x"5e",
    x"3e",
    x"06",
    x"cd",
    x"93",
    x"00",
    x"18",
    x"07",
    x"3a",
    x"8c",
    x"e1",
    x"a7",
    x"c4",
    x"08",
    x"90",
    x"21",
    x"90",
    x"e1",
    x"06",
    x"01",
    x"cd",
    x"e1",
    x"8a",
    x"21",
    x"90",
    x"e1",
    x"11",
    x"98",
    x"91",
    x"0e",
    x"03",
    x"06",
    x"29",
    x"d5",
    x"e5",
    x"7e",
    x"a7",
    x"c4",
    x"b1",
    x"90",
    x"e1",
    x"11",
    x"08",
    x"00",
    x"19",
    x"d1",
    x"13",
    x"13",
    x"10",
    x"ef",
    x"c9",
    x"3d",
    x"c2",
    x"c4",
    x"90",
    x"e5",
    x"34",
    x"23",
    x"23",
    x"36",
    x"fe",
    x"23",
    x"23",
    x"1a",
    x"77",
    x"13",
    x"23",
    x"1a",
    x"77",
    x"e1",
    x"23",
    x"56",
    x"23",
    x"34",
    x"7e",
    x"ba",
    x"da",
    x"4a",
    x"91",
    x"36",
    x"00",
    x"23",
    x"23",
    x"5e",
    x"23",
    x"56",
    x"1a",
    x"13",
    x"fe",
    x"d0",
    x"da",
    x"3d",
    x"91",
    x"fe",
    x"f0",
    x"38",
    x"31",
    x"e5",
    x"21",
    x"e8",
    x"90",
    x"e6",
    x"0f",
    x"c3",
    x"f8",
    x"8a",
    x"f4",
    x"90",
    x"07",
    x"91",
    x"1b",
    x"91",
    x"25",
    x"91",
    x"2d",
    x"91",
    x"35",
    x"91",
    x"e1",
    x"23",
    x"13",
    x"13",
    x"73",
    x"23",
    x"72",
    x"2b",
    x"2b",
    x"1b",
    x"1a",
    x"1b",
    x"08",
    x"1a",
    x"5f",
    x"08",
    x"57",
    x"18",
    x"cd",
    x"e1",
    x"23",
    x"5e",
    x"23",
    x"56",
    x"2b",
    x"2b",
    x"18",
    x"c4",
    x"e5",
    x"2b",
    x"2b",
    x"2b",
    x"2b",
    x"d6",
    x"d0",
    x"77",
    x"e1",
    x"18",
    x"b9",
    x"e1",
    x"2b",
    x"2b",
    x"1a",
    x"13",
    x"77",
    x"23",
    x"23",
    x"18",
    x"af",
    x"e1",
    x"2b",
    x"2b",
    x"34",
    x"23",
    x"23",
    x"18",
    x"a7",
    x"e1",
    x"2b",
    x"2b",
    x"35",
    x"23",
    x"23",
    x"18",
    x"9f",
    x"e1",
    x"11",
    x"fb",
    x"ff",
    x"19",
    x"36",
    x"00",
    x"c9",
    x"72",
    x"2b",
    x"73",
    x"2b",
    x"7e",
    x"e6",
    x"60",
    x"28",
    x"03",
    x"32",
    x"8c",
    x"e1",
    x"2b",
    x"0d",
    x"f8",
    x"23",
    x"7e",
    x"08",
    x"23",
    x"5e",
    x"23",
    x"56",
    x"1b",
    x"1a",
    x"e6",
    x"f0",
    x"fe",
    x"e0",
    x"28",
    x"38",
    x"21",
    x"ea",
    x"91",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"cb",
    x"3f",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"1a",
    x"e6",
    x"0f",
    x"cb",
    x"3c",
    x"cb",
    x"1d",
    x"3d",
    x"20",
    x"f9",
    x"eb",
    x"79",
    x"87",
    x"87",
    x"21",
    x"80",
    x"e1",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"73",
    x"23",
    x"72",
    x"23",
    x"08",
    x"57",
    x"e6",
    x"1f",
    x"77",
    x"23",
    x"af",
    x"cb",
    x"12",
    x"17",
    x"77",
    x"c9",
    x"21",
    x"00",
    x"00",
    x"18",
    x"df",
    x"d1",
    x"8f",
    x"ee",
    x"8f",
    x"f4",
    x"8f",
    x"ad",
    x"8f",
    x"b9",
    x"8f",
    x"91",
    x"8f",
    x"9f",
    x"8f",
    x"f4",
    x"8f",
    x"02",
    x"92",
    x"30",
    x"95",
    x"1b",
    x"8f",
    x"3e",
    x"8f",
    x"53",
    x"8f",
    x"82",
    x"8f",
    x"a9",
    x"93",
    x"27",
    x"94",
    x"c5",
    x"8f",
    x"14",
    x"92",
    x"4b",
    x"92",
    x"54",
    x"95",
    x"78",
    x"95",
    x"23",
    x"92",
    x"5a",
    x"92",
    x"82",
    x"92",
    x"b8",
    x"92",
    x"fb",
    x"92",
    x"3e",
    x"93",
    x"82",
    x"93",
    x"8f",
    x"93",
    x"9c",
    x"93",
    x"53",
    x"94",
    x"5c",
    x"94",
    x"02",
    x"95",
    x"ba",
    x"94",
    x"b8",
    x"92",
    x"b0",
    x"92",
    x"fa",
    x"8f",
    x"a6",
    x"92",
    x"b5",
    x"93",
    x"e2",
    x"93",
    x"11",
    x"94",
    x"c8",
    x"d5",
    x"c8",
    x"c9",
    x"75",
    x"be",
    x"c4",
    x"b3",
    x"ad",
    x"a9",
    x"28",
    x"a0",
    x"2a",
    x"97",
    x"ae",
    x"8e",
    x"ac",
    x"86",
    x"1d",
    x"7f",
    x"fb",
    x"77",
    x"3f",
    x"71",
    x"f2",
    x"50",
    x"da",
    x"97",
    x"b7",
    x"08",
    x"b7",
    x"97",
    x"87",
    x"67",
    x"87",
    x"97",
    x"57",
    x"47",
    x"07",
    x"97",
    x"97",
    x"f5",
    x"d5",
    x"f0",
    x"38",
    x"92",
    x"96",
    x"b6",
    x"07",
    x"27",
    x"07",
    x"47",
    x"67",
    x"87",
    x"e4",
    x"97",
    x"f5",
    x"d6",
    x"f0",
    x"38",
    x"92",
    x"96",
    x"07",
    x"b6",
    x"27",
    x"07",
    x"47",
    x"27",
    x"57",
    x"47",
    x"97",
    x"87",
    x"97",
    x"b7",
    x"47",
    x"67",
    x"87",
    x"f5",
    x"f2",
    x"50",
    x"48",
    x"08",
    x"28",
    x"b7",
    x"08",
    x"97",
    x"b7",
    x"87",
    x"97",
    x"47",
    x"57",
    x"27",
    x"07",
    x"b6",
    x"96",
    x"86",
    x"f1",
    x"d5",
    x"f0",
    x"6f",
    x"92",
    x"46",
    x"56",
    x"66",
    x"86",
    x"96",
    x"b6",
    x"07",
    x"27",
    x"e4",
    x"47",
    x"f5",
    x"d6",
    x"f0",
    x"6f",
    x"92",
    x"46",
    x"86",
    x"66",
    x"96",
    x"86",
    x"07",
    x"b6",
    x"27",
    x"07",
    x"47",
    x"27",
    x"57",
    x"47",
    x"27",
    x"07",
    x"b6",
    x"f5",
    x"f2",
    x"0d",
    x"08",
    x"97",
    x"b7",
    x"87",
    x"97",
    x"67",
    x"87",
    x"47",
    x"57",
    x"07",
    x"27",
    x"b6",
    x"96",
    x"86",
    x"66",
    x"46",
    x"f1",
    x"d6",
    x"f2",
    x"0d",
    x"95",
    x"95",
    x"46",
    x"46",
    x"96",
    x"96",
    x"96",
    x"46",
    x"26",
    x"06",
    x"b5",
    x"95",
    x"95",
    x"b5",
    x"b5",
    x"b5",
    x"06",
    x"06",
    x"26",
    x"26",
    x"46",
    x"46",
    x"56",
    x"56",
    x"46",
    x"46",
    x"26",
    x"06",
    x"b5",
    x"85",
    x"95",
    x"b5",
    x"f5",
    x"f2",
    x"0b",
    x"d6",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"f0",
    x"bb",
    x"92",
    x"f2",
    x"0d",
    x"d6",
    x"c0",
    x"c0",
    x"f0",
    x"bb",
    x"92",
    x"f2",
    x"0f",
    x"d6",
    x"77",
    x"77",
    x"77",
    x"08",
    x"28",
    x"28",
    x"28",
    x"58",
    x"48",
    x"48",
    x"48",
    x"08",
    x"28",
    x"28",
    x"28",
    x"98",
    x"78",
    x"78",
    x"78",
    x"08",
    x"28",
    x"28",
    x"28",
    x"58",
    x"48",
    x"48",
    x"48",
    x"08",
    x"78",
    x"78",
    x"78",
    x"b8",
    x"09",
    x"09",
    x"09",
    x"a8",
    x"88",
    x"88",
    x"88",
    x"78",
    x"58",
    x"58",
    x"58",
    x"38",
    x"28",
    x"28",
    x"28",
    x"a7",
    x"a8",
    x"a8",
    x"a8",
    x"09",
    x"a8",
    x"a8",
    x"a8",
    x"78",
    x"d8",
    x"98",
    x"58",
    x"28",
    x"78",
    x"48",
    x"28",
    x"f5",
    x"f2",
    x"0d",
    x"d6",
    x"48",
    x"48",
    x"48",
    x"77",
    x"28",
    x"28",
    x"28",
    x"97",
    x"08",
    x"08",
    x"08",
    x"77",
    x"97",
    x"97",
    x"97",
    x"b7",
    x"48",
    x"48",
    x"48",
    x"77",
    x"28",
    x"28",
    x"28",
    x"97",
    x"08",
    x"08",
    x"08",
    x"77",
    x"28",
    x"28",
    x"28",
    x"78",
    x"88",
    x"88",
    x"88",
    x"78",
    x"58",
    x"58",
    x"58",
    x"38",
    x"28",
    x"28",
    x"28",
    x"08",
    x"a7",
    x"a7",
    x"a7",
    x"28",
    x"38",
    x"38",
    x"38",
    x"58",
    x"38",
    x"38",
    x"38",
    x"08",
    x"d8",
    x"58",
    x"28",
    x"97",
    x"28",
    x"b7",
    x"97",
    x"f5",
    x"f2",
    x"0d",
    x"d6",
    x"77",
    x"77",
    x"77",
    x"77",
    x"97",
    x"97",
    x"97",
    x"08",
    x"b7",
    x"b7",
    x"b7",
    x"b7",
    x"77",
    x"77",
    x"77",
    x"77",
    x"08",
    x"08",
    x"08",
    x"08",
    x"28",
    x"28",
    x"28",
    x"58",
    x"48",
    x"48",
    x"48",
    x"48",
    x"28",
    x"28",
    x"28",
    x"28",
    x"38",
    x"38",
    x"38",
    x"38",
    x"28",
    x"28",
    x"28",
    x"08",
    x"a7",
    x"a7",
    x"a7",
    x"a7",
    x"38",
    x"38",
    x"38",
    x"38",
    x"a8",
    x"a8",
    x"a8",
    x"a8",
    x"78",
    x"78",
    x"78",
    x"38",
    x"28",
    x"28",
    x"28",
    x"28",
    x"78",
    x"78",
    x"78",
    x"48",
    x"f5",
    x"f2",
    x"0d",
    x"d7",
    x"28",
    x"28",
    x"c0",
    x"28",
    x"38",
    x"58",
    x"78",
    x"78",
    x"78",
    x"f5",
    x"f2",
    x"0d",
    x"d7",
    x"97",
    x"97",
    x"c0",
    x"97",
    x"a7",
    x"08",
    x"28",
    x"28",
    x"28",
    x"f5",
    x"f2",
    x"0d",
    x"d7",
    x"67",
    x"67",
    x"c0",
    x"67",
    x"77",
    x"97",
    x"b7",
    x"b7",
    x"b7",
    x"f5",
    x"f2",
    x"0f",
    x"d4",
    x"77",
    x"97",
    x"77",
    x"97",
    x"08",
    x"28",
    x"08",
    x"28",
    x"f5",
    x"e8",
    x"f2",
    x"50",
    x"b7",
    x"77",
    x"47",
    x"07",
    x"e2",
    x"c0",
    x"d6",
    x"b7",
    x"e2",
    x"77",
    x"d6",
    x"47",
    x"d8",
    x"07",
    x"47",
    x"77",
    x"37",
    x"67",
    x"97",
    x"e8",
    x"57",
    x"97",
    x"08",
    x"28",
    x"e2",
    x"c0",
    x"d6",
    x"38",
    x"e2",
    x"08",
    x"d6",
    x"87",
    x"d8",
    x"57",
    x"37",
    x"07",
    x"87",
    x"37",
    x"08",
    x"f0",
    x"b5",
    x"93",
    x"e8",
    x"f2",
    x"10",
    x"77",
    x"47",
    x"07",
    x"b6",
    x"d6",
    x"c0",
    x"c0",
    x"c0",
    x"76",
    x"47",
    x"47",
    x"47",
    x"07",
    x"d8",
    x"b6",
    x"07",
    x"47",
    x"07",
    x"37",
    x"57",
    x"e8",
    x"27",
    x"57",
    x"97",
    x"08",
    x"d6",
    x"c0",
    x"c0",
    x"c0",
    x"08",
    x"87",
    x"87",
    x"87",
    x"57",
    x"d8",
    x"37",
    x"07",
    x"86",
    x"57",
    x"37",
    x"86",
    x"f0",
    x"e2",
    x"93",
    x"f2",
    x"0d",
    x"e8",
    x"b7",
    x"b7",
    x"b7",
    x"b7",
    x"b7",
    x"b7",
    x"77",
    x"b7",
    x"97",
    x"97",
    x"97",
    x"97",
    x"87",
    x"87",
    x"08",
    x"28",
    x"f0",
    x"11",
    x"94",
    x"f2",
    x"0e",
    x"d3",
    x"0a",
    x"b9",
    x"a9",
    x"99",
    x"89",
    x"79",
    x"69",
    x"59",
    x"49",
    x"39",
    x"29",
    x"19",
    x"09",
    x"b8",
    x"a8",
    x"98",
    x"88",
    x"78",
    x"68",
    x"58",
    x"48",
    x"38",
    x"28",
    x"18",
    x"08",
    x"b7",
    x"a7",
    x"97",
    x"87",
    x"77",
    x"67",
    x"57",
    x"47",
    x"37",
    x"27",
    x"17",
    x"07",
    x"b6",
    x"a6",
    x"96",
    x"f5",
    x"f2",
    x"0f",
    x"d1",
    x"b8",
    x"c0",
    x"78",
    x"c0",
    x"98",
    x"f5",
    x"d5",
    x"f2",
    x"4f",
    x"48",
    x"48",
    x"f3",
    x"48",
    x"48",
    x"f4",
    x"48",
    x"f3",
    x"48",
    x"f4",
    x"28",
    x"28",
    x"28",
    x"f3",
    x"28",
    x"f4",
    x"28",
    x"28",
    x"28",
    x"f3",
    x"28",
    x"f4",
    x"28",
    x"f3",
    x"28",
    x"d5",
    x"f4",
    x"58",
    x"58",
    x"f3",
    x"58",
    x"58",
    x"f4",
    x"58",
    x"f3",
    x"58",
    x"f4",
    x"48",
    x"48",
    x"48",
    x"f3",
    x"48",
    x"f4",
    x"48",
    x"48",
    x"48",
    x"f3",
    x"48",
    x"f4",
    x"48",
    x"f3",
    x"48",
    x"58",
    x"58",
    x"c0",
    x"58",
    x"f4",
    x"58",
    x"f3",
    x"58",
    x"78",
    x"78",
    x"c0",
    x"78",
    x"f4",
    x"78",
    x"f3",
    x"78",
    x"f4",
    x"78",
    x"f3",
    x"78",
    x"f4",
    x"78",
    x"f3",
    x"78",
    x"98",
    x"98",
    x"c0",
    x"98",
    x"f4",
    x"98",
    x"f3",
    x"98",
    x"f4",
    x"98",
    x"f3",
    x"98",
    x"f0",
    x"27",
    x"94",
    x"f2",
    x"0e",
    x"d5",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"07",
    x"47",
    x"77",
    x"08",
    x"f2",
    x"10",
    x"18",
    x"18",
    x"c0",
    x"18",
    x"f4",
    x"18",
    x"f3",
    x"18",
    x"38",
    x"38",
    x"c0",
    x"38",
    x"f4",
    x"38",
    x"f3",
    x"38",
    x"f4",
    x"38",
    x"f3",
    x"38",
    x"f4",
    x"38",
    x"f3",
    x"38",
    x"f2",
    x"0d",
    x"57",
    x"97",
    x"08",
    x"58",
    x"58",
    x"08",
    x"97",
    x"57",
    x"f5",
    x"f2",
    x"0d",
    x"e4",
    x"07",
    x"76",
    x"07",
    x"76",
    x"07",
    x"76",
    x"07",
    x"76",
    x"d5",
    x"f2",
    x"10",
    x"86",
    x"86",
    x"c0",
    x"86",
    x"f4",
    x"86",
    x"f3",
    x"86",
    x"a6",
    x"a6",
    x"c0",
    x"a6",
    x"f4",
    x"a6",
    x"f3",
    x"a6",
    x"f4",
    x"a6",
    x"f3",
    x"a6",
    x"f4",
    x"a6",
    x"f3",
    x"a6",
    x"f2",
    x"0f",
    x"da",
    x"58",
    x"58",
    x"08",
    x"57",
    x"f5",
    x"f2",
    x"50",
    x"d6",
    x"48",
    x"18",
    x"28",
    x"b7",
    x"08",
    x"97",
    x"b7",
    x"87",
    x"97",
    x"47",
    x"67",
    x"27",
    x"17",
    x"b6",
    x"96",
    x"86",
    x"96",
    x"17",
    x"b6",
    x"27",
    x"17",
    x"47",
    x"27",
    x"67",
    x"47",
    x"97",
    x"87",
    x"97",
    x"b7",
    x"47",
    x"67",
    x"87",
    x"f5",
    x"f2",
    x"0d",
    x"d6",
    x"18",
    x"97",
    x"b7",
    x"87",
    x"97",
    x"67",
    x"87",
    x"47",
    x"67",
    x"17",
    x"27",
    x"b6",
    x"96",
    x"86",
    x"66",
    x"46",
    x"46",
    x"96",
    x"86",
    x"b6",
    x"96",
    x"17",
    x"b6",
    x"27",
    x"17",
    x"47",
    x"27",
    x"67",
    x"47",
    x"27",
    x"17",
    x"b6",
    x"f5",
    x"f2",
    x"0d",
    x"d6",
    x"95",
    x"95",
    x"46",
    x"46",
    x"96",
    x"96",
    x"96",
    x"46",
    x"26",
    x"16",
    x"b5",
    x"95",
    x"95",
    x"b5",
    x"b5",
    x"b5",
    x"16",
    x"16",
    x"26",
    x"26",
    x"46",
    x"46",
    x"66",
    x"66",
    x"46",
    x"46",
    x"26",
    x"16",
    x"b5",
    x"85",
    x"95",
    x"b5",
    x"f5",
    x"fd",
    x"21",
    x"0c",
    x"98",
    x"fd",
    x"7e",
    x"00",
    x"fd",
    x"23",
    x"a7",
    x"ca",
    x"ae",
    x"98",
    x"47",
    x"e6",
    x"3f",
    x"cb",
    x"78",
    x"28",
    x"08",
    x"21",
    x"fd",
    x"95",
    x"cd",
    x"f8",
    x"8a",
    x"18",
    x"e8",
    x"cb",
    x"70",
    x"28",
    x"05",
    x"cd",
    x"17",
    x"96",
    x"18",
    x"df",
    x"cd",
    x"28",
    x"96",
    x"18",
    x"da",
    x"87",
    x"21",
    x"ed",
    x"95",
    x"85",
    x"6f",
    x"30",
    x"01",
    x"24",
    x"7e",
    x"23",
    x"66",
    x"6f",
    x"7e",
    x"32",
    x"5c",
    x"e0",
    x"23",
    x"e5",
    x"dd",
    x"e1",
    x"11",
    x"00",
    x"f0",
    x"cd",
    x"33",
    x"96",
    x"11",
    x"00",
    x"3c",
    x"21",
    x"00",
    x"f0",
    x"01",
    x"00",
    x"01",
    x"c3",
    x"5c",
    x"00",
    x"4d",
    x"9e",
    x"8f",
    x"9e",
    x"c0",
    x"9e",
    x"f1",
    x"9e",
    x"22",
    x"9f",
    x"64",
    x"9d",
    x"23",
    x"9d",
    x"53",
    x"9f",
    x"33",
    x"96",
    x"80",
    x"96",
    x"b7",
    x"96",
    x"c3",
    x"96",
    x"f0",
    x"96",
    x"d9",
    x"96",
    x"32",
    x"97",
    x"46",
    x"97",
    x"5e",
    x"97",
    x"65",
    x"97",
    x"75",
    x"97",
    x"84",
    x"97",
    x"06",
    x"97",
    x"06",
    x"00",
    x"87",
    x"87",
    x"87",
    x"cb",
    x"10",
    x"4f",
    x"dd",
    x"e5",
    x"e1",
    x"ed",
    x"b0",
    x"e5",
    x"dd",
    x"e1",
    x"c9",
    x"26",
    x"00",
    x"87",
    x"87",
    x"87",
    x"cb",
    x"14",
    x"6f",
    x"19",
    x"eb",
    x"c9",
    x"3e",
    x"02",
    x"cd",
    x"17",
    x"96",
    x"dd",
    x"7e",
    x"00",
    x"3c",
    x"20",
    x"09",
    x"dd",
    x"23",
    x"3e",
    x"06",
    x"cd",
    x"17",
    x"96",
    x"18",
    x"08",
    x"cd",
    x"d9",
    x"96",
    x"3e",
    x"04",
    x"cd",
    x"17",
    x"96",
    x"dd",
    x"7e",
    x"00",
    x"3c",
    x"20",
    x"09",
    x"21",
    x"00",
    x"f0",
    x"01",
    x"c0",
    x"00",
    x"ed",
    x"b0",
    x"c9",
    x"cd",
    x"64",
    x"96",
    x"cd",
    x"64",
    x"96",
    x"cd",
    x"67",
    x"96",
    x"21",
    x"c8",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"d0",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"b0",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"b8",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"c9",
    x"3e",
    x"01",
    x"cd",
    x"17",
    x"96",
    x"21",
    x"08",
    x"00",
    x"19",
    x"d5",
    x"eb",
    x"21",
    x"f0",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"f8",
    x"ff",
    x"cd",
    x"a4",
    x"96",
    x"d1",
    x"21",
    x"10",
    x"00",
    x"cd",
    x"a4",
    x"96",
    x"21",
    x"10",
    x"00",
    x"19",
    x"eb",
    x"c9",
    x"19",
    x"0e",
    x"08",
    x"06",
    x"08",
    x"e5",
    x"cb",
    x"06",
    x"1f",
    x"23",
    x"10",
    x"fa",
    x"e1",
    x"12",
    x"13",
    x"0d",
    x"20",
    x"f1",
    x"c9",
    x"3e",
    x"01",
    x"cd",
    x"28",
    x"96",
    x"3e",
    x"02",
    x"cd",
    x"17",
    x"96",
    x"18",
    x"05",
    x"3e",
    x"03",
    x"cd",
    x"17",
    x"96",
    x"21",
    x"f8",
    x"ff",
    x"cd",
    x"f5",
    x"96",
    x"21",
    x"e8",
    x"ff",
    x"cd",
    x"f5",
    x"96",
    x"21",
    x"d8",
    x"ff",
    x"18",
    x"1c",
    x"21",
    x"f0",
    x"ff",
    x"e5",
    x"cd",
    x"e1",
    x"96",
    x"e1",
    x"cd",
    x"f5",
    x"96",
    x"21",
    x"f8",
    x"ff",
    x"19",
    x"06",
    x"08",
    x"cb",
    x"26",
    x"23",
    x"10",
    x"fb",
    x"c9",
    x"21",
    x"f8",
    x"ff",
    x"18",
    x"ec",
    x"19",
    x"0e",
    x"08",
    x"06",
    x"08",
    x"cb",
    x"06",
    x"1f",
    x"10",
    x"fb",
    x"12",
    x"23",
    x"13",
    x"0d",
    x"20",
    x"f3",
    x"c9",
    x"cd",
    x"12",
    x"97",
    x"cd",
    x"0f",
    x"97",
    x"cd",
    x"0f",
    x"97",
    x"cd",
    x"12",
    x"97",
    x"d5",
    x"21",
    x"d0",
    x"ff",
    x"19",
    x"01",
    x"30",
    x"00",
    x"ed",
    x"b0",
    x"e1",
    x"0e",
    x"06",
    x"af",
    x"08",
    x"af",
    x"06",
    x"08",
    x"08",
    x"cb",
    x"1f",
    x"cb",
    x"1e",
    x"23",
    x"10",
    x"f9",
    x"cb",
    x"1f",
    x"0d",
    x"20",
    x"f1",
    x"c9",
    x"3e",
    x"01",
    x"cd",
    x"17",
    x"96",
    x"3e",
    x"01",
    x"cd",
    x"28",
    x"96",
    x"3e",
    x"01",
    x"cd",
    x"17",
    x"96",
    x"3e",
    x"01",
    x"c3",
    x"28",
    x"96",
    x"3e",
    x"01",
    x"cd",
    x"17",
    x"96",
    x"3e",
    x"01",
    x"cd",
    x"28",
    x"96",
    x"21",
    x"e0",
    x"ff",
    x"19",
    x"01",
    x"08",
    x"00",
    x"ed",
    x"b0",
    x"3e",
    x"01",
    x"c3",
    x"28",
    x"96",
    x"cd",
    x"6a",
    x"97",
    x"e5",
    x"dd",
    x"e1",
    x"c9",
    x"cd",
    x"6a",
    x"97",
    x"eb",
    x"c9",
    x"fd",
    x"6e",
    x"00",
    x"fd",
    x"23",
    x"fd",
    x"66",
    x"00",
    x"fd",
    x"23",
    x"c9",
    x"d5",
    x"cd",
    x"65",
    x"97",
    x"21",
    x"00",
    x"e8",
    x"01",
    x"00",
    x"08",
    x"cd",
    x"5c",
    x"00",
    x"d1",
    x"c9",
    x"21",
    x"00",
    x"f3",
    x"06",
    x"b0",
    x"cd",
    x"e1",
    x"8a",
    x"11",
    x"00",
    x"e8",
    x"c9",
    x"dd",
    x"21",
    x"ec",
    x"97",
    x"11",
    x"00",
    x"f0",
    x"06",
    x"03",
    x"c5",
    x"dd",
    x"6e",
    x"00",
    x"dd",
    x"23",
    x"dd",
    x"66",
    x"00",
    x"dd",
    x"23",
    x"cd",
    x"c2",
    x"97",
    x"c1",
    x"10",
    x"ef",
    x"11",
    x"00",
    x"05",
    x"21",
    x"00",
    x"f0",
    x"01",
    x"80",
    x"01",
    x"cd",
    x"5c",
    x"00",
    x"11",
    x"00",
    x"1c",
    x"21",
    x"f2",
    x"97",
    x"01",
    x"1a",
    x"00",
    x"c3",
    x"5c",
    x"00",
    x"06",
    x"04",
    x"c5",
    x"46",
    x"23",
    x"4e",
    x"23",
    x"3e",
    x"08",
    x"08",
    x"78",
    x"41",
    x"4f",
    x"af",
    x"cb",
    x"11",
    x"30",
    x"02",
    x"f6",
    x"f0",
    x"cb",
    x"11",
    x"30",
    x"02",
    x"f6",
    x"0f",
    x"12",
    x"13",
    x"12",
    x"13",
    x"12",
    x"13",
    x"12",
    x"13",
    x"08",
    x"3d",
    x"20",
    x"e3",
    x"c1",
    x"10",
    x"d9",
    x"c9",
    x"53",
    x"9a",
    x"23",
    x"9a",
    x"7b",
    x"9a",
    x"60",
    x"60",
    x"60",
    x"60",
    x"60",
    x"60",
    x"f0",
    x"f0",
    x"f0",
    x"f0",
    x"f0",
    x"f0",
    x"70",
    x"70",
    x"70",
    x"70",
    x"70",
    x"70",
    x"c0",
    x"40",
    x"40",
    x"40",
    x"40",
    x"40",
    x"40",
    x"40",
    x"8b",
    x"88",
    x"1b",
    x"9a",
    x"60",
    x"08",
    x"88",
    x"7b",
    x"99",
    x"54",
    x"04",
    x"60",
    x"88",
    x"bb",
    x"99",
    x"4c",
    x"04",
    x"60",
    x"88",
    x"d3",
    x"9c",
    x"42",
    x"85",
    x"42",
    x"85",
    x"88",
    x"d3",
    x"9c",
    x"42",
    x"85",
    x"42",
    x"85",
    x"8a",
    x"00",
    x"00",
    x"89",
    x"80",
    x"ec",
    x"88",
    x"1b",
    x"9b",
    x"41",
    x"84",
    x"41",
    x"84",
    x"04",
    x"83",
    x"8a",
    x"00",
    x"08",
    x"89",
    x"80",
    x"ec",
    x"83",
    x"83",
    x"83",
    x"83",
    x"83",
    x"83",
    x"45",
    x"84",
    x"41",
    x"84",
    x"41",
    x"84",
    x"41",
    x"84",
    x"45",
    x"84",
    x"41",
    x"84",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"81",
    x"8a",
    x"00",
    x"10",
    x"8b",
    x"88",
    x"a3",
    x"9c",
    x"80",
    x"88",
    x"e3",
    x"9c",
    x"80",
    x"88",
    x"24",
    x"9d",
    x"80",
    x"88",
    x"65",
    x"9d",
    x"80",
    x"20",
    x"81",
    x"81",
    x"81",
    x"81",
    x"80",
    x"44",
    x"86",
    x"87",
    x"87",
    x"87",
    x"87",
    x"86",
    x"87",
    x"8a",
    x"00",
    x"38",
    x"8b",
    x"89",
    x"00",
    x"e9",
    x"88",
    x"24",
    x"9d",
    x"42",
    x"85",
    x"02",
    x"8c",
    x"89",
    x"80",
    x"ea",
    x"88",
    x"13",
    x"9d",
    x"42",
    x"85",
    x"02",
    x"8c",
    x"89",
    x"00",
    x"ec",
    x"88",
    x"65",
    x"9d",
    x"42",
    x"85",
    x"02",
    x"8c",
    x"89",
    x"80",
    x"ed",
    x"88",
    x"54",
    x"9d",
    x"42",
    x"85",
    x"02",
    x"8c",
    x"00",
    x"11",
    x"e6",
    x"98",
    x"21",
    x"00",
    x"20",
    x"1a",
    x"13",
    x"a7",
    x"c8",
    x"47",
    x"cb",
    x"7f",
    x"28",
    x"10",
    x"e6",
    x"70",
    x"c6",
    x"10",
    x"e5",
    x"6f",
    x"26",
    x"00",
    x"78",
    x"29",
    x"29",
    x"44",
    x"4d",
    x"e1",
    x"18",
    x"0b",
    x"e6",
    x"70",
    x"0f",
    x"0f",
    x"0f",
    x"0f",
    x"3c",
    x"4f",
    x"78",
    x"06",
    x"00",
    x"e6",
    x"0f",
    x"07",
    x"07",
    x"07",
    x"07",
    x"c5",
    x"cd",
    x"56",
    x"00",
    x"c1",
    x"09",
    x"18",
    x"ce",
    x"d6",
    x"df",
    x"d7",
    x"84",
    x"8c",
    x"d9",
    x"d9",
    x"ba",
    x"96",
    x"df",
    x"d7",
    x"8f",
    x"76",
    x"57",
    x"66",
    x"27",
    x"46",
    x"27",
    x"57",
    x"16",
    x"76",
    x"76",
    x"76",
    x"d5",
    x"d5",
    x"ba",
    x"96",
    x"df",
    x"da",
    x"7f",
    x"34",
    x"17",
    x"36",
    x"24",
    x"27",
    x"16",
    x"24",
    x"27",
    x"34",
    x"17",
    x"16",
    x"7f",
    x"76",
    x"06",
    x"24",
    x"27",
    x"36",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"06",
    x"24",
    x"27",
    x"06",
    x"7f",
    x"24",
    x"27",
    x"26",
    x"24",
    x"27",
    x"36",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"06",
    x"24",
    x"27",
    x"06",
    x"24",
    x"27",
    x"16",
    x"24",
    x"17",
    x"36",
    x"24",
    x"27",
    x"36",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"06",
    x"24",
    x"27",
    x"06",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"36",
    x"24",
    x"27",
    x"36",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"06",
    x"24",
    x"27",
    x"06",
    x"24",
    x"27",
    x"16",
    x"24",
    x"47",
    x"06",
    x"24",
    x"37",
    x"26",
    x"24",
    x"17",
    x"26",
    x"24",
    x"17",
    x"16",
    x"14",
    x"37",
    x"24",
    x"47",
    x"7b",
    x"7b",
    x"79",
    x"79",
    x"74",
    x"74",
    x"74",
    x"74",
    x"7d",
    x"7d",
    x"7d",
    x"7d",
    x"7a",
    x"7a",
    x"7a",
    x"7a",
    x"7c",
    x"7c",
    x"7c",
    x"7c",
    x"ef",
    x"00",
    x"3f",
    x"3f",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"8f",
    x"cf",
    x"c0",
    x"cf",
    x"df",
    x"d8",
    x"df",
    x"cf",
    x"cf",
    x"ef",
    x"6c",
    x"ec",
    x"ec",
    x"6c",
    x"ec",
    x"ec",
    x"f8",
    x"fd",
    x"cd",
    x"cd",
    x"cd",
    x"cd",
    x"cd",
    x"cc",
    x"fe",
    x"fe",
    x"80",
    x"80",
    x"80",
    x"80",
    x"fe",
    x"fe",
    x"7e",
    x"ff",
    x"c3",
    x"c3",
    x"c3",
    x"c3",
    x"ff",
    x"7e",
    x"7f",
    x"7f",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"80",
    x"80",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"1c",
    x"26",
    x"63",
    x"63",
    x"63",
    x"32",
    x"1c",
    x"00",
    x"0c",
    x"1c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"3f",
    x"00",
    x"3e",
    x"63",
    x"07",
    x"1e",
    x"3c",
    x"70",
    x"7f",
    x"00",
    x"3f",
    x"06",
    x"0c",
    x"1e",
    x"03",
    x"63",
    x"3e",
    x"00",
    x"0e",
    x"1e",
    x"36",
    x"66",
    x"7f",
    x"06",
    x"06",
    x"00",
    x"7e",
    x"60",
    x"7e",
    x"03",
    x"03",
    x"63",
    x"3e",
    x"00",
    x"1c",
    x"30",
    x"60",
    x"7e",
    x"61",
    x"61",
    x"3e",
    x"00",
    x"7f",
    x"63",
    x"06",
    x"0c",
    x"18",
    x"18",
    x"18",
    x"00",
    x"3c",
    x"62",
    x"72",
    x"3c",
    x"4f",
    x"43",
    x"3e",
    x"00",
    x"3e",
    x"63",
    x"63",
    x"3f",
    x"03",
    x"06",
    x"3c",
    x"00",
    x"60",
    x"78",
    x"7e",
    x"78",
    x"60",
    x"60",
    x"60",
    x"00",
    x"21",
    x"52",
    x"24",
    x"08",
    x"12",
    x"25",
    x"42",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"1c",
    x"36",
    x"63",
    x"63",
    x"7f",
    x"63",
    x"63",
    x"00",
    x"7e",
    x"63",
    x"63",
    x"7e",
    x"63",
    x"63",
    x"7e",
    x"00",
    x"1e",
    x"33",
    x"60",
    x"60",
    x"60",
    x"33",
    x"1e",
    x"00",
    x"7c",
    x"66",
    x"63",
    x"63",
    x"63",
    x"66",
    x"7c",
    x"00",
    x"3f",
    x"30",
    x"30",
    x"3e",
    x"30",
    x"30",
    x"3f",
    x"00",
    x"7f",
    x"60",
    x"60",
    x"7e",
    x"60",
    x"60",
    x"60",
    x"00",
    x"1f",
    x"30",
    x"60",
    x"67",
    x"63",
    x"33",
    x"1f",
    x"00",
    x"63",
    x"63",
    x"63",
    x"7f",
    x"63",
    x"63",
    x"63",
    x"00",
    x"3f",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"3f",
    x"00",
    x"03",
    x"03",
    x"03",
    x"03",
    x"03",
    x"63",
    x"3e",
    x"00",
    x"63",
    x"66",
    x"6c",
    x"78",
    x"7c",
    x"6e",
    x"67",
    x"00",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"3f",
    x"00",
    x"63",
    x"77",
    x"7f",
    x"7f",
    x"6b",
    x"63",
    x"63",
    x"00",
    x"63",
    x"73",
    x"7b",
    x"7f",
    x"6f",
    x"67",
    x"63",
    x"00",
    x"3e",
    x"63",
    x"63",
    x"63",
    x"63",
    x"63",
    x"3e",
    x"00",
    x"7e",
    x"63",
    x"63",
    x"63",
    x"7e",
    x"60",
    x"60",
    x"00",
    x"3e",
    x"63",
    x"63",
    x"63",
    x"6f",
    x"66",
    x"3d",
    x"00",
    x"7e",
    x"63",
    x"63",
    x"67",
    x"7c",
    x"6e",
    x"67",
    x"00",
    x"3c",
    x"66",
    x"60",
    x"3e",
    x"03",
    x"63",
    x"3e",
    x"00",
    x"3f",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"00",
    x"63",
    x"63",
    x"63",
    x"63",
    x"63",
    x"63",
    x"3e",
    x"00",
    x"63",
    x"63",
    x"63",
    x"77",
    x"3e",
    x"1c",
    x"08",
    x"00",
    x"63",
    x"63",
    x"6b",
    x"7f",
    x"7f",
    x"77",
    x"63",
    x"00",
    x"63",
    x"77",
    x"3e",
    x"1c",
    x"3e",
    x"77",
    x"63",
    x"00",
    x"33",
    x"33",
    x"33",
    x"1e",
    x"0c",
    x"0c",
    x"0c",
    x"00",
    x"7f",
    x"07",
    x"0e",
    x"1c",
    x"38",
    x"70",
    x"7f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"3c",
    x"3c",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"7f",
    x"7f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"18",
    x"18",
    x"00",
    x"18",
    x"3c",
    x"3c",
    x"18",
    x"18",
    x"00",
    x"18",
    x"00",
    x"3c",
    x"42",
    x"9d",
    x"a1",
    x"a1",
    x"9d",
    x"42",
    x"3c",
    x"01",
    x"01",
    x"01",
    x"03",
    x"03",
    x"13",
    x"13",
    x"17",
    x"9e",
    x"9c",
    x"bd",
    x"ff",
    x"ff",
    x"ef",
    x"cd",
    x"81",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"01",
    x"00",
    x"00",
    x"03",
    x"20",
    x"20",
    x"10",
    x"0c",
    x"03",
    x"c0",
    x"38",
    x"07",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"04",
    x"03",
    x"00",
    x"08",
    x"07",
    x"00",
    x"0e",
    x"e0",
    x"1f",
    x"80",
    x"70",
    x"0f",
    x"00",
    x"f0",
    x"0f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"18",
    x"07",
    x"00",
    x"30",
    x"0e",
    x"01",
    x"70",
    x"e0",
    x"1f",
    x"00",
    x"f0",
    x"0f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"0f",
    x"c0",
    x"3c",
    x"03",
    x"00",
    x"f0",
    x"0f",
    x"e0",
    x"c0",
    x"3f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"c0",
    x"3f",
    x"02",
    x"01",
    x"00",
    x"04",
    x"03",
    x"00",
    x"07",
    x"00",
    x"1f",
    x"c0",
    x"3c",
    x"03",
    x"80",
    x"78",
    x"07",
    x"f0",
    x"80",
    x"7f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"c0",
    x"3f",
    x"08",
    x"07",
    x"00",
    x"10",
    x"0f",
    x"00",
    x"3e",
    x"01",
    x"0f",
    x"80",
    x"78",
    x"07",
    x"00",
    x"f0",
    x"0f",
    x"e0",
    x"80",
    x"7f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"c0",
    x"3f",
    x"70",
    x"0f",
    x"00",
    x"60",
    x"1e",
    x"01",
    x"00",
    x"00",
    x"1f",
    x"00",
    x"f0",
    x"0f",
    x"00",
    x"e0",
    x"1f",
    x"00",
    x"80",
    x"7f",
    x"00",
    x"c0",
    x"3f",
    x"00",
    x"80",
    x"7f",
    x"00",
    x"00",
    x"00",
    x"00",
    x"fe",
    x"fe",
    x"00",
    x"fe",
    x"fe",
    x"00",
    x"fe",
    x"ba",
    x"d6",
    x"6c",
    x"38",
    x"10",
    x"00",
    x"00",
    x"fe",
    x"00",
    x"7c",
    x"60",
    x"7c",
    x"0c",
    x"7c",
    x"00",
    x"fe",
    x"fe",
    x"ba",
    x"54",
    x"28",
    x"10",
    x"00",
    x"00",
    x"7f",
    x"7e",
    x"7c",
    x"46",
    x"72",
    x"60",
    x"78",
    x"72",
    x"3a",
    x"1a",
    x"0e",
    x"07",
    x"03",
    x"01",
    x"ff",
    x"fe",
    x"fc",
    x"e6",
    x"c2",
    x"98",
    x"bc",
    x"9e",
    x"ce",
    x"67",
    x"30",
    x"1b",
    x"08",
    x"07",
    x"03",
    x"01",
    x"ff",
    x"fc",
    x"dc",
    x"8c",
    x"80",
    x"90",
    x"84",
    x"80",
    x"fe",
    x"7e",
    x"96",
    x"62",
    x"02",
    x"12",
    x"42",
    x"02",
    x"aa",
    x"3c",
    x"3c",
    x"18",
    x"0b",
    x"07",
    x"03",
    x"01",
    x"aa",
    x"78",
    x"78",
    x"30",
    x"a0",
    x"c0",
    x"80",
    x"00",
    x"ff",
    x"ff",
    x"c3",
    x"c3",
    x"ff",
    x"c3",
    x"c3",
    x"ff",
    x"e1",
    x"70",
    x"38",
    x"1c",
    x"0e",
    x"07",
    x"03",
    x"01",
    x"00",
    x"00",
    x"60",
    x"10",
    x"0c",
    x"05",
    x"02",
    x"0c",
    x"00",
    x"11",
    x"67",
    x"0e",
    x"1d",
    x"1b",
    x"1b",
    x"0d",
    x"00",
    x"00",
    x"00",
    x"1b",
    x"3f",
    x"3a",
    x"6a",
    x"77",
    x"be",
    x"dd",
    x"d2",
    x"94",
    x"c9",
    x"a2",
    x"88",
    x"d2",
    x"80",
    x"40",
    x"28",
    x"10",
    x"67",
    x"0f",
    x"1a",
    x"1d",
    x"1e",
    x"c7",
    x"22",
    x"ae",
    x"6d",
    x"2e",
    x"1d",
    x"3a",
    x"1e",
    x"3f",
    x"35",
    x"1a",
    x"b5",
    x"ea",
    x"55",
    x"aa",
    x"a8",
    x"5a",
    x"2d",
    x"da",
    x"22",
    x"49",
    x"25",
    x"4a",
    x"00",
    x"00",
    x"20",
    x"12",
    x"09",
    x"05",
    x"02",
    x"0c",
    x"01",
    x"03",
    x"86",
    x"6d",
    x"2d",
    x"66",
    x"2f",
    x"0d",
    x"08",
    x"08",
    x"24",
    x"40",
    x"1f",
    x"3e",
    x"39",
    x"5f",
    x"d2",
    x"14",
    x"2b",
    x"89",
    x"54",
    x"29",
    x"e4",
    x"12",
    x"01",
    x"01",
    x"01",
    x"03",
    x"03",
    x"13",
    x"13",
    x"17",
    x"9e",
    x"9c",
    x"bd",
    x"ff",
    x"ff",
    x"ef",
    x"cd",
    x"81",
    x"00",
    x"00",
    x"00",
    x"09",
    x"12",
    x"26",
    x"7f",
    x"fe",
    x"1f",
    x"1f",
    x"07",
    x"0b",
    x"13",
    x"00",
    x"00",
    x"00",
    x"00",
    x"02",
    x"04",
    x"18",
    x"38",
    x"70",
    x"e0",
    x"40",
    x"48",
    x"f0",
    x"e0",
    x"c8",
    x"d0",
    x"e0",
    x"c0",
    x"80",
    x"02",
    x"02",
    x"1f",
    x"09",
    x"07",
    x"19",
    x"38",
    x"f8",
    x"75",
    x"32",
    x"32",
    x"38",
    x"18",
    x"0c",
    x"06",
    x"02",
    x"02",
    x"02",
    x"1f",
    x"09",
    x"07",
    x"09",
    x"38",
    x"f8",
    x"7d",
    x"5a",
    x"d2",
    x"b0",
    x"90",
    x"90",
    x"f0",
    x"60",
    x"00",
    x"08",
    x"0e",
    x"3e",
    x"77",
    x"ce",
    x"b9",
    x"f3",
    x"e4",
    x"c0",
    x"01",
    x"00",
    x"00",
    x"01",
    x"03",
    x"03",
    x"20",
    x"34",
    x"6a",
    x"ec",
    x"32",
    x"3f",
    x"0c",
    x"88",
    x"d8",
    x"bc",
    x"3c",
    x"6e",
    x"d8",
    x"d8",
    x"30",
    x"e0",
    x"00",
    x"00",
    x"00",
    x"12",
    x"32",
    x"35",
    x"37",
    x"3f",
    x"0c",
    x"1f",
    x"3e",
    x"3b",
    x"19",
    x"00",
    x"00",
    x"00",
    x"09",
    x"00",
    x"00",
    x"00",
    x"12",
    x"72",
    x"75",
    x"77",
    x"3f",
    x"1c",
    x"3f",
    x"7e",
    x"3b",
    x"08",
    x"00",
    x"00",
    x"00",
    x"00",
    x"06",
    x"0f",
    x"0e",
    x"0c",
    x"7d",
    x"7f",
    x"7d",
    x"3e",
    x"2d",
    x"0f",
    x"07",
    x"01",
    x"03",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"20",
    x"c0",
    x"48",
    x"f0",
    x"d0",
    x"e4",
    x"4e",
    x"fe",
    x"fc",
    x"e0",
    x"e0",
    x"e0",
    x"00",
    x"00",
    x"00",
    x"00",
    x"11",
    x"17",
    x"0d",
    x"07",
    x"0c",
    x"0f",
    x"1a",
    x"3a",
    x"3b",
    x"39",
    x"00",
    x"00",
    x"00",
    x"05",
    x"00",
    x"00",
    x"00",
    x"21",
    x"17",
    x"0d",
    x"07",
    x"0c",
    x"1f",
    x"3a",
    x"7a",
    x"73",
    x"71",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"01",
    x"01",
    x"00",
    x"7d",
    x"ff",
    x"fa",
    x"67",
    x"0d",
    x"0b",
    x"0e",
    x"00",
    x"01",
    x"01",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"d0",
    x"60",
    x"f0",
    x"50",
    x"6e",
    x"c0",
    x"60",
    x"e0",
    x"e0",
    x"e0",
    x"e0",
    x"c0",
    x"00",
    x"06",
    x"2c",
    x"20",
    x"5b",
    x"52",
    x"05",
    x"65",
    x"00",
    x"02",
    x"1d",
    x"25",
    x"56",
    x"49",
    x"1e",
    x"25",
    x"00",
    x"66",
    x"89",
    x"63",
    x"2c",
    x"c5",
    x"ba",
    x"25",
    x"00",
    x"32",
    x"6d",
    x"09",
    x"64",
    x"18",
    x"a3",
    x"94",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"01",
    x"03",
    x"03",
    x"01",
    x"01",
    x"01",
    x"01",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"01",
    x"02",
    x"04",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"10",
    x"e0",
    x"e0",
    x"e0",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"40",
    x"40",
    x"e0",
    x"e0",
    x"40",
    x"40",
    x"40",
    x"40",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"02",
    x"02",
    x"07",
    x"07",
    x"02",
    x"02",
    x"02",
    x"02",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"08",
    x"19",
    x"29",
    x"49",
    x"7d",
    x"09",
    x"08",
    x"00",
    x"c6",
    x"29",
    x"29",
    x"29",
    x"29",
    x"29",
    x"c6",
    x"00",
    x"38",
    x"45",
    x"45",
    x"39",
    x"45",
    x"45",
    x"38",
    x"00",
    x"98",
    x"a5",
    x"a5",
    x"a5",
    x"a5",
    x"a5",
    x"98",
    x"00",
    x"bc",
    x"a1",
    x"a1",
    x"b9",
    x"85",
    x"85",
    x"b8",
    x"00",
    x"98",
    x"a1",
    x"a1",
    x"b9",
    x"a5",
    x"a5",
    x"98",
    x"00",
    x"62",
    x"95",
    x"15",
    x"25",
    x"45",
    x"85",
    x"f2",
    x"00",
    x"22",
    x"55",
    x"55",
    x"55",
    x"55",
    x"55",
    x"22",
    x"00",
    x"f2",
    x"15",
    x"65",
    x"15",
    x"15",
    x"95",
    x"62",
    x"0d",
    x"00",
    x"00",
    x"00",
    x"02",
    x"2a",
    x"39",
    x"1b",
    x"1b",
    x"07",
    x"03",
    x"03",
    x"11",
    x"09",
    x"06",
    x"00",
    x"00",
    x"ff",
    x"00",
    x"00",
    x"00",
    x"80",
    x"a8",
    x"38",
    x"b0",
    x"b0",
    x"e0",
    x"80",
    x"80",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"02",
    x"03",
    x"07",
    x"06",
    x"05",
    x"03",
    x"07",
    x"07",
    x"07",
    x"08",
    x"08",
    x"07",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"80",
    x"20",
    x"50",
    x"e0",
    x"c8",
    x"d8",
    x"bc",
    x"70",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"03",
    x"00",
    x"00",
    x"01",
    x"01",
    x"05",
    x"0d",
    x"03",
    x"1f",
    x"1f",
    x"3f",
    x"33",
    x"21",
    x"21",
    x"01",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"0e",
    x"1f",
    x"2f",
    x"03",
    x"03",
    x"03",
    x"04",
    x"08",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"c8",
    x"50",
    x"20",
    x"d8",
    x"c8",
    x"e0",
    x"f0",
    x"70",
    x"70",
    x"20",
    x"40",
    x"00",
    x"00",
    x"0a",
    x"00",
    x"00",
    x"00",
    x"01",
    x"23",
    x"27",
    x"3f",
    x"2b",
    x"37",
    x"1d",
    x"0d",
    x"05",
    x"01",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"06",
    x"0c",
    x"1c",
    x"17",
    x"13",
    x"1f",
    x"1f",
    x"13",
    x"05",
    x"09",
    x"13",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"e0",
    x"e0",
    x"e0",
    x"e0",
    x"e4",
    x"bc",
    x"98",
    x"f0",
    x"00",
    x"00",
    x"00",
    x"07",
    x"00",
    x"00",
    x"06",
    x"02",
    x"01",
    x"fd",
    x"7f",
    x"1d",
    x"01",
    x"01",
    x"01",
    x"01",
    x"01",
    x"00",
    x"00",
    x"00",
    x"04",
    x"06",
    x"0f",
    x"0f",
    x"07",
    x"07",
    x"03",
    x"00",
    x"01",
    x"02",
    x"04",
    x"08",
    x"10",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"10",
    x"30",
    x"9c",
    x"a8",
    x"c0",
    x"f0",
    x"7c",
    x"7e",
    x"3f",
    x"0c",
    x"00",
    x"00",
    x"00",
    x"00",
    x"04",
    x"06",
    x"0e",
    x"1f",
    x"1c",
    x"19",
    x"1c",
    x"5f",
    x"6f",
    x"67",
    x"71",
    x"7b",
    x"7f",
    x"6f",
    x"67",
    x"03",
    x"03",
    x"00",
    x"04",
    x"0d",
    x"1d",
    x"39",
    x"7d",
    x"f9",
    x"d8",
    x"1f",
    x"1f",
    x"0f",
    x"1f",
    x"3b",
    x"30",
    x"00",
    x"00",
    x"7c",
    x"fc",
    x"fb",
    x"87",
    x"97",
    x"c7",
    x"e7",
    x"fe",
    x"7c",
    x"00",
    x"2e",
    x"fc",
    x"f8",
    x"70",
    x"e0",
    x"c0",
    x"06",
    x"80",
    x"50",
    x"20",
    x"50",
    x"08",
    x"05",
    x"03",
    x"03",
    x"1f",
    x"7f",
    x"7d",
    x"f1",
    x"c3",
    x"03",
    x"03",
    x"02",
    x"ff",
    x"20",
    x"60",
    x"e0",
    x"e0",
    x"c2",
    x"de",
    x"fc",
    x"f8",
    x"30",
    x"90",
    x"f8",
    x"bc",
    x"8c",
    x"00",
    x"00",
    x"00",
    x"80",
    x"50",
    x"20",
    x"50",
    x"08",
    x"06",
    x"7f",
    x"ff",
    x"ff",
    x"3f",
    x"03",
    x"03",
    x"03",
    x"03",
    x"03",
    x"02",
    x"10",
    x"30",
    x"70",
    x"70",
    x"f0",
    x"e0",
    x"e0",
    x"c0",
    x"38",
    x"9e",
    x"fe",
    x"fc",
    x"8c",
    x"00",
    x"00",
    x"00",
    x"ff",
    x"42",
    x"59",
    x"20",
    x"46",
    x"55",
    x"4b",
    x"41",
    x"53",
    x"48",
    x"49",
    x"e4",
    x"e5",
    x"e8",
    x"ec",
    x"ec",
    x"f2",
    x"f9",
    x"00",
    x"00",
    x"07",
    x"0e",
    x"14",
    x"14",
    x"18",
    x"1b",
    x"1c",
    x"1c",
    x"1b",
    x"18",
    x"14",
    x"14",
    x"0e",
    x"07",
    x"00",
    x"00",
    x"f9",
    x"f2",
    x"ec",
    x"ec",
    x"e8",
    x"e5",
    x"e4",
    x"d8",
    x"d9",
    x"dd",
    x"e4",
    x"e4",
    x"ec",
    x"f6",
    x"00",
    x"00",
    x"0a",
    x"14",
    x"1c",
    x"1c",
    x"23",
    x"27",
    x"28",
    x"28",
    x"27",
    x"23",
    x"1c",
    x"1c",
    x"14",
    x"0a",
    x"00",
    x"00",
    x"f6",
    x"ec",
    x"e4",
    x"e4",
    x"dd",
    x"d9",
    x"d8",
    x"c8",
    x"ca",
    x"d0",
    x"d8",
    x"d8",
    x"e4",
    x"f2",
    x"00",
    x"00",
    x"0e",
    x"1c",
    x"28",
    x"28",
    x"30",
    x"36",
    x"38",
    x"38",
    x"36",
    x"30",
    x"28",
    x"28",
    x"1c",
    x"0e",
    x"00",
    x"00",
    x"f2",
    x"e4",
    x"d8",
    x"d8",
    x"d0",
    x"ca",
    x"c8"
);
begin

process (cs)
begin
if rising_edge(cs) then
    D <= galaga(to_integer(unsigned(A)));
end if;
end process;
end;

